

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  INV_X1 U322 ( .A(n560), .ZN(n540) );
  XNOR2_X2 U323 ( .A(KEYINPUT126), .B(n456), .ZN(n566) );
  NOR2_X1 U324 ( .A1(n578), .A2(n365), .ZN(n366) );
  XNOR2_X1 U325 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U326 ( .A(n481), .B(n480), .ZN(n505) );
  XNOR2_X1 U327 ( .A(n325), .B(n324), .ZN(n529) );
  XOR2_X1 U328 ( .A(G78GAT), .B(G148GAT), .Z(n290) );
  XNOR2_X1 U329 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n470) );
  XNOR2_X1 U330 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U331 ( .A(KEYINPUT85), .ZN(n315) );
  INV_X1 U332 ( .A(KEYINPUT78), .ZN(n354) );
  XNOR2_X1 U333 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U336 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U337 ( .A(n440), .B(n294), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n357), .B(n356), .ZN(n360) );
  XOR2_X1 U339 ( .A(n578), .B(KEYINPUT41), .Z(n553) );
  XNOR2_X1 U340 ( .A(n305), .B(n304), .ZN(n578) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n482) );
  XNOR2_X1 U342 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U343 ( .A(n482), .B(KEYINPUT40), .ZN(n483) );
  XNOR2_X1 U344 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XNOR2_X1 U345 ( .A(n484), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G85GAT), .B(G57GAT), .Z(n416) );
  XOR2_X1 U347 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n329) );
  XOR2_X1 U348 ( .A(n416), .B(n329), .Z(n305) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n291) );
  XNOR2_X1 U350 ( .A(n290), .B(n291), .ZN(n440) );
  NAND2_X1 U351 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  INV_X1 U352 ( .A(KEYINPUT70), .ZN(n292) );
  XOR2_X1 U353 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n296) );
  XNOR2_X1 U354 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n295) );
  XOR2_X1 U355 ( .A(n296), .B(n295), .Z(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n303) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n299), .B(G120GAT), .ZN(n318) );
  XOR2_X1 U359 ( .A(G64GAT), .B(G92GAT), .Z(n301) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n396) );
  XNOR2_X1 U362 ( .A(n318), .B(n396), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U364 ( .A(KEYINPUT109), .B(n553), .ZN(n533) );
  INV_X1 U365 ( .A(n533), .ZN(n457) );
  XOR2_X1 U366 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n307) );
  XNOR2_X1 U367 ( .A(G190GAT), .B(KEYINPUT64), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U369 ( .A(G176GAT), .B(KEYINPUT83), .Z(n309) );
  XNOR2_X1 U370 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U372 ( .A(n311), .B(n310), .Z(n321) );
  XOR2_X1 U373 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n313) );
  XNOR2_X1 U374 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U375 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U376 ( .A(G169GAT), .B(n314), .Z(n397) );
  NAND2_X1 U377 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n397), .B(n319), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n323) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n322), .B(KEYINPUT80), .ZN(n417) );
  XOR2_X1 U382 ( .A(n323), .B(n417), .Z(n325) );
  XOR2_X1 U383 ( .A(G43GAT), .B(G134GAT), .Z(n348) );
  XOR2_X1 U384 ( .A(G15GAT), .B(G127GAT), .Z(n328) );
  XNOR2_X1 U385 ( .A(n348), .B(n328), .ZN(n324) );
  XOR2_X1 U386 ( .A(G155GAT), .B(G78GAT), .Z(n327) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G211GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n342) );
  XOR2_X1 U389 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U392 ( .A(G64GAT), .B(KEYINPUT15), .Z(n333) );
  XNOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U396 ( .A(G1GAT), .B(G8GAT), .Z(n373) );
  XOR2_X1 U397 ( .A(KEYINPUT14), .B(G57GAT), .Z(n337) );
  XNOR2_X1 U398 ( .A(G183GAT), .B(G71GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n373), .B(n338), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n536) );
  INV_X1 U403 ( .A(n536), .ZN(n581) );
  XOR2_X1 U404 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n344) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n352) );
  XOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n346) );
  XNOR2_X1 U408 ( .A(G218GAT), .B(KEYINPUT75), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U410 ( .A(n347), .B(G92GAT), .Z(n350) );
  XNOR2_X1 U411 ( .A(G99GAT), .B(n348), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U413 ( .A(n352), .B(n351), .Z(n362) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n353), .B(KEYINPUT77), .ZN(n400) );
  XOR2_X1 U416 ( .A(G50GAT), .B(G162GAT), .Z(n446) );
  XNOR2_X1 U417 ( .A(n400), .B(n446), .ZN(n357) );
  AND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n358), .B(KEYINPUT8), .ZN(n377) );
  XNOR2_X1 U421 ( .A(n377), .B(KEYINPUT9), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n560) );
  XOR2_X1 U424 ( .A(KEYINPUT36), .B(n540), .Z(n583) );
  NAND2_X1 U425 ( .A1(n581), .A2(n583), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n363), .B(KEYINPUT117), .ZN(n364) );
  XOR2_X1 U427 ( .A(KEYINPUT45), .B(n364), .Z(n365) );
  XNOR2_X1 U428 ( .A(KEYINPUT118), .B(n366), .ZN(n385) );
  XOR2_X1 U429 ( .A(KEYINPUT29), .B(G113GAT), .Z(n368) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G15GAT), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U432 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n370) );
  XNOR2_X1 U433 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U436 ( .A(G197GAT), .B(G43GAT), .Z(n375) );
  XOR2_X1 U437 ( .A(G141GAT), .B(G22GAT), .Z(n447) );
  XNOR2_X1 U438 ( .A(n447), .B(n373), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n376), .B(G36GAT), .Z(n382) );
  XOR2_X1 U441 ( .A(n377), .B(KEYINPUT68), .Z(n379) );
  NAND2_X1 U442 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n380), .B(G50GAT), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U446 ( .A(n384), .B(n383), .Z(n549) );
  NAND2_X1 U447 ( .A1(n385), .A2(n549), .ZN(n394) );
  XOR2_X1 U448 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n386) );
  XNOR2_X1 U449 ( .A(KEYINPUT114), .B(n386), .ZN(n388) );
  INV_X1 U450 ( .A(n549), .ZN(n574) );
  NAND2_X1 U451 ( .A1(n574), .A2(n553), .ZN(n387) );
  XOR2_X1 U452 ( .A(n388), .B(n387), .Z(n389) );
  NOR2_X1 U453 ( .A1(n581), .A2(n389), .ZN(n390) );
  NAND2_X1 U454 ( .A1(n390), .A2(n540), .ZN(n392) );
  XOR2_X1 U455 ( .A(KEYINPUT116), .B(KEYINPUT47), .Z(n391) );
  NAND2_X1 U456 ( .A1(n394), .A2(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(KEYINPUT48), .B(n395), .Z(n546) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n399) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U462 ( .A(n401), .B(n400), .Z(n405) );
  XOR2_X1 U463 ( .A(G211GAT), .B(KEYINPUT21), .Z(n403) );
  XNOR2_X1 U464 ( .A(G197GAT), .B(G218GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n441) );
  XNOR2_X1 U466 ( .A(G8GAT), .B(n441), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n520) );
  XOR2_X1 U469 ( .A(n520), .B(KEYINPUT125), .Z(n408) );
  NOR2_X1 U470 ( .A1(n546), .A2(n408), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n409), .B(KEYINPUT54), .ZN(n571) );
  XOR2_X1 U472 ( .A(G148GAT), .B(G127GAT), .Z(n411) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U475 ( .A(KEYINPUT76), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(G134GAT), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n434) );
  XOR2_X1 U479 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U482 ( .A(n420), .B(KEYINPUT1), .Z(n424) );
  XOR2_X1 U483 ( .A(G155GAT), .B(KEYINPUT3), .Z(n422) );
  XNOR2_X1 U484 ( .A(KEYINPUT89), .B(KEYINPUT2), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n444) );
  XNOR2_X1 U486 ( .A(n444), .B(KEYINPUT91), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U488 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n426) );
  XNOR2_X1 U489 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n425) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U491 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n428) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n427) );
  XNOR2_X1 U493 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U494 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n570) );
  XOR2_X1 U497 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U500 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n438) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U503 ( .A(n439), .B(G204GAT), .Z(n443) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U506 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n469) );
  INV_X1 U510 ( .A(n469), .ZN(n452) );
  AND2_X1 U511 ( .A1(n570), .A2(n452), .ZN(n453) );
  AND2_X1 U512 ( .A1(n571), .A2(n453), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n529), .A2(n455), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n457), .A2(n566), .ZN(n460) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n481) );
  OR2_X1 U518 ( .A1(n578), .A2(n549), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT73), .ZN(n488) );
  XNOR2_X1 U520 ( .A(n529), .B(KEYINPUT86), .ZN(n463) );
  XOR2_X1 U521 ( .A(n520), .B(KEYINPUT27), .Z(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT28), .B(n469), .Z(n526) );
  NAND2_X1 U523 ( .A1(n466), .A2(n526), .ZN(n462) );
  NOR2_X1 U524 ( .A1(n570), .A2(n462), .ZN(n531) );
  NAND2_X1 U525 ( .A1(n463), .A2(n531), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(KEYINPUT98), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n469), .A2(n529), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT26), .ZN(n573) );
  INV_X1 U529 ( .A(n466), .ZN(n467) );
  NOR2_X1 U530 ( .A1(n573), .A2(n467), .ZN(n548) );
  NOR2_X1 U531 ( .A1(n529), .A2(n520), .ZN(n468) );
  NOR2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n471) );
  NOR2_X1 U533 ( .A1(n548), .A2(n472), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(n473), .Z(n474) );
  NAND2_X1 U535 ( .A1(n474), .A2(n570), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(n477), .ZN(n487) );
  NOR2_X1 U538 ( .A1(n581), .A2(n487), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n583), .A2(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n479), .ZN(n518) );
  NAND2_X1 U541 ( .A1(n488), .A2(n518), .ZN(n480) );
  NOR2_X1 U542 ( .A1(n529), .A2(n505), .ZN(n484) );
  NAND2_X1 U543 ( .A1(n540), .A2(n581), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(n485), .ZN(n486) );
  NOR2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n507) );
  NAND2_X1 U546 ( .A1(n507), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(KEYINPUT102), .ZN(n498) );
  NOR2_X1 U548 ( .A1(n498), .A2(n570), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT103), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n498), .A2(n520), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(n493), .Z(n494) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n494), .ZN(G1325GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n496) );
  NOR2_X1 U556 ( .A1(n529), .A2(n498), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n497), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n498), .A2(n526), .ZN(n499) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n499), .Z(G1327GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n501) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT108), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U564 ( .A1(n505), .A2(n570), .ZN(n502) );
  XOR2_X1 U565 ( .A(n503), .B(n502), .Z(G1328GAT) );
  NOR2_X1 U566 ( .A1(n505), .A2(n520), .ZN(n504) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n505), .A2(n526), .ZN(n506) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  NOR2_X1 U570 ( .A1(n574), .A2(n533), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n507), .A2(n517), .ZN(n513) );
  NOR2_X1 U572 ( .A1(n570), .A2(n513), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n520), .A2(n513), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n529), .A2(n513), .ZN(n512) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n570), .A2(n525), .ZN(n519) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n525), .ZN(n521) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n529), .A2(n525), .ZN(n522) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n524) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT113), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U595 ( .A(n528), .B(n527), .Z(G1339GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n546), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n541) );
  NOR2_X1 U598 ( .A1(n549), .A2(n541), .ZN(n532) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n541), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n541), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n543) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT121), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n570), .A2(n546), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n552) );
  NOR2_X1 U614 ( .A1(n549), .A2(n552), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(n550), .Z(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT124), .Z(n555) );
  INV_X1 U618 ( .A(n552), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(n556), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n561), .A2(n581), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  BUF_X1 U626 ( .A(n560), .Z(n565) );
  NAND2_X1 U627 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n566), .A2(n574), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n581), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n584), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

