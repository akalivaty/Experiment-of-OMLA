//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n204), .A2(KEYINPUT71), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT71), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n203), .C1(new_n206), .C2(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  AND2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT74), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT74), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n226), .B2(G141gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n216), .B1(new_n228), .B2(new_n217), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n215), .B(new_n220), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n214), .B1(new_n231), .B2(KEYINPUT29), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n228), .ZN(new_n233));
  INV_X1    g032(.A(new_n216), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n223), .B2(new_n225), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n237), .B2(new_n222), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n220), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n232), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(KEYINPUT81), .B(new_n239), .C1(new_n240), .C2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g047(.A(new_n222), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT74), .B(G148gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(new_n236), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n236), .A2(G148gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n228), .B1(new_n222), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n251), .A2(new_n235), .B1(new_n253), .B2(new_n218), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT29), .B1(new_n254), .B2(new_n215), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT82), .B1(new_n255), .B2(new_n213), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n214), .B(new_n257), .C1(new_n231), .C2(KEYINPUT29), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n247), .A2(new_n248), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n245), .B1(new_n259), .B2(new_n242), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261));
  OAI21_X1  g060(.A(G22gat), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g061(.A(KEYINPUT84), .B(new_n245), .C1(new_n259), .C2(new_n242), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n202), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n242), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n244), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT84), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n261), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(KEYINPUT85), .A3(G22gat), .A4(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT83), .B(G22gat), .Z(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G50gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G78gat), .B(G106gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n264), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n275), .B(KEYINPUT80), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n266), .A2(new_n270), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n271), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n277), .A2(KEYINPUT86), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT86), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AND4_X1   g099(.A1(new_n287), .A2(new_n294), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT66), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT23), .B(new_n296), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n286), .A2(new_n298), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n311), .A2(new_n290), .A3(new_n293), .A4(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(new_n307), .A3(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n301), .A2(new_n303), .B1(new_n314), .B2(new_n299), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n285), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n298), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n320), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n318), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n319), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n315), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT72), .B(new_n284), .C1(new_n330), .C2(KEYINPUT29), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n299), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n286), .A2(new_n298), .A3(new_n299), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n303), .A2(new_n334), .A3(new_n294), .A4(new_n295), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n327), .A3(new_n328), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT29), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n284), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n315), .B2(new_n329), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(KEYINPUT73), .A3(new_n337), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n331), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n214), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n339), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n214), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n214), .B2(new_n345), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(KEYINPUT30), .A3(new_n359), .ZN(new_n360));
  OR3_X1    g159(.A1(new_n352), .A2(KEYINPUT30), .A3(new_n355), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n364), .B1(KEYINPUT1), .B2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G113gat), .B(G120gat), .Z(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n315), .B2(new_n329), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n366), .A2(new_n370), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n336), .A2(new_n373), .A3(new_n337), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n363), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT32), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n375), .A2(KEYINPUT33), .ZN(new_n378));
  XOR2_X1   g177(.A(G15gat), .B(G43gat), .Z(new_n379));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n375), .B2(KEYINPUT33), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n363), .A3(new_n374), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT34), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT34), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n382), .A2(new_n386), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n389), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n383), .A2(new_n385), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n383), .A2(new_n385), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n373), .A2(new_n402), .A3(new_n254), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT4), .B1(new_n239), .B2(new_n371), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n254), .A2(new_n215), .B1(new_n370), .B2(new_n366), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT75), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n230), .A2(new_n371), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n215), .B1(new_n238), .B2(new_n220), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n401), .B(new_n405), .C1(new_n408), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n373), .A2(new_n254), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n239), .A2(new_n371), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n401), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n407), .A2(KEYINPUT75), .A3(new_n230), .A4(new_n371), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n419), .A2(new_n420), .B1(new_n404), .B2(new_n403), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n418), .B1(new_n421), .B2(new_n401), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  INV_X1    g223(.A(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT0), .B(G57gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT6), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n415), .B(new_n428), .C1(new_n422), .C2(new_n414), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n362), .A2(new_n399), .A3(new_n400), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n283), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n277), .A2(new_n280), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n277), .A2(KEYINPUT86), .A3(new_n280), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n444));
  INV_X1    g243(.A(new_n418), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n413), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n428), .A4(new_n415), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n414), .B1(new_n413), .B2(new_n445), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT5), .B1(new_n421), .B2(new_n401), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n429), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n454), .B2(new_n433), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n451), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n434), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n362), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT78), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n444), .B(new_n449), .C1(new_n430), .C2(new_n451), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n430), .A2(new_n451), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n435), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n362), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT69), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n443), .A2(new_n460), .A3(new_n465), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n438), .B1(new_n470), .B2(KEYINPUT35), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n443), .B1(new_n460), .B2(new_n465), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT70), .B(KEYINPUT36), .C1(new_n393), .C2(new_n397), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n398), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n346), .A2(new_n351), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n355), .B1(new_n357), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT90), .B(new_n355), .C1(new_n357), .C2(new_n482), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n357), .A2(new_n480), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n345), .A2(new_n213), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n348), .A2(new_n349), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n490), .B2(new_n214), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n488), .A2(new_n492), .A3(new_n479), .A4(new_n355), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n432), .A3(new_n435), .A4(new_n359), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n405), .B1(new_n408), .B2(new_n412), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  INV_X1    g295(.A(new_n401), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n416), .A2(new_n417), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n496), .B1(new_n499), .B2(new_n401), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n421), .B2(new_n401), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n501), .A3(new_n429), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT40), .B1(new_n502), .B2(KEYINPUT87), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n501), .A3(new_n504), .A4(new_n429), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n431), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n360), .A2(new_n361), .A3(new_n514), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n487), .A2(new_n494), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n478), .B1(new_n283), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n472), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n471), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G15gat), .B(G22gat), .Z(new_n520));
  INV_X1    g319(.A(G1gat), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT91), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(G8gat), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528));
  NAND2_X1  g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  NOR2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(KEYINPUT94), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n526), .B1(new_n537), .B2(KEYINPUT21), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n537), .A2(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT95), .ZN(new_n545));
  XOR2_X1   g344(.A(G183gat), .B(G211gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n543), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(new_n550), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT101), .B(G92gat), .Z(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT100), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n558), .B2(KEYINPUT100), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n557), .A2(new_n425), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT99), .B(new_n563), .C1(new_n425), .C2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT99), .B1(new_n425), .B2(new_n564), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G99gat), .B(G106gat), .Z(new_n571));
  AOI21_X1  g370(.A(new_n556), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n570), .B(new_n571), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n556), .ZN(new_n574));
  OR3_X1    g373(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n575), .A2(new_n576), .B1(G29gat), .B2(G36gat), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n578));
  XNOR2_X1  g377(.A(G43gat), .B(G50gat), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n577), .A2(KEYINPUT15), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(KEYINPUT17), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(new_n589), .A3(new_n582), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n573), .A2(new_n556), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n588), .B(new_n590), .C1(new_n591), .C2(new_n572), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n555), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  AND4_X1   g392(.A1(new_n555), .A2(new_n592), .A3(new_n585), .A4(new_n586), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT98), .ZN(new_n597));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  OAI21_X1  g398(.A(KEYINPUT103), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601));
  INV_X1    g400(.A(new_n599), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n601), .B(new_n602), .C1(new_n593), .C2(new_n594), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n593), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n605), .B2(KEYINPUT104), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(KEYINPUT104), .B2(new_n595), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n526), .A2(new_n584), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n525), .A3(new_n590), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n612), .A2(KEYINPUT92), .B1(G229gat), .B2(G233gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(KEYINPUT92), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n525), .B(new_n583), .ZN(new_n617));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  AOI22_X1  g418(.A1(new_n614), .A2(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n610), .A2(new_n611), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n615), .A3(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G197gat), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT11), .B(G169gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n622), .A3(new_n628), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n623), .A2(KEYINPUT93), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G230gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n537), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n574), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n573), .A2(new_n537), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n537), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n636), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n639), .B1(new_n574), .B2(new_n637), .ZN(new_n645));
  INV_X1    g444(.A(new_n636), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G204gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(G176gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n644), .A2(new_n647), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n635), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR4_X1   g457(.A1(new_n519), .A2(new_n554), .A3(new_n609), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n458), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n459), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT16), .B(G8gat), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT106), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(G8gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(G1325gat));
  AOI21_X1  g467(.A(G15gat), .B1(new_n659), .B2(new_n399), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n478), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n478), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n669), .B1(new_n659), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n283), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n460), .A2(new_n465), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n469), .B1(new_n281), .B2(new_n282), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT35), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n438), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n463), .A2(new_n464), .A3(new_n362), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n464), .B1(new_n463), .B2(new_n362), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n283), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n485), .A2(new_n486), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT38), .ZN(new_n689));
  INV_X1    g488(.A(new_n494), .ZN(new_n690));
  INV_X1    g489(.A(new_n509), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT88), .B1(new_n503), .B2(new_n505), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n360), .A2(new_n361), .A3(new_n514), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n689), .A2(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n443), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n687), .A2(new_n696), .A3(new_n478), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n684), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n553), .A2(new_n658), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n609), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n463), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n608), .A2(KEYINPUT44), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n471), .A2(new_n518), .A3(KEYINPUT109), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n684), .B2(new_n697), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n519), .B2(new_n608), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n704), .B1(new_n711), .B2(new_n699), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n705), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT109), .B1(new_n471), .B2(new_n518), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n685), .A2(new_n686), .ZN(new_n716));
  INV_X1    g515(.A(new_n681), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n400), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n707), .B(new_n697), .C1(new_n718), .C2(new_n438), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n714), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n698), .B2(new_n609), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n704), .B(new_n699), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n463), .B1(new_n713), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(G29gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n703), .B1(new_n724), .B2(new_n725), .ZN(G1328gat));
  NOR2_X1   g525(.A1(new_n519), .A2(new_n608), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n362), .A2(G36gat), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n727), .A2(new_n728), .A3(new_n699), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n729), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT111), .B1(new_n700), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n362), .B1(new_n713), .B2(new_n723), .ZN(new_n738));
  INV_X1    g537(.A(G36gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(G1329gat));
  NAND2_X1  g539(.A1(new_n711), .A2(new_n699), .ZN(new_n741));
  OAI21_X1  g540(.A(G43gat), .B1(new_n741), .B2(new_n478), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n700), .A2(G43gat), .A3(new_n398), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n723), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n674), .B1(new_n712), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n743), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  OR2_X1    g548(.A1(new_n700), .A2(KEYINPUT114), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n443), .A2(G50gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n700), .A2(KEYINPUT114), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n750), .A2(new_n756), .A3(new_n753), .A4(new_n751), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G50gat), .B1(new_n741), .B2(new_n443), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT48), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n752), .A2(new_n754), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n283), .B1(new_n712), .B2(new_n746), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n715), .A2(new_n719), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n458), .B(KEYINPUT116), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n553), .A2(new_n608), .A3(new_n635), .ZN(new_n768));
  INV_X1    g567(.A(new_n656), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  OAI21_X1  g571(.A(new_n770), .B1(new_n706), .B2(new_n708), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT117), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n766), .A2(new_n775), .A3(new_n770), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n362), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n773), .B2(new_n398), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n774), .A2(new_n776), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n673), .A2(new_n782), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n775), .B1(new_n766), .B2(new_n770), .ZN(new_n788));
  INV_X1    g587(.A(new_n770), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT117), .B(new_n789), .C1(new_n715), .C2(new_n719), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n784), .B(new_n786), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n783), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n783), .B(new_n795), .C1(new_n787), .C2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n785), .A2(new_n283), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT119), .B(G78gat), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1335gat));
  INV_X1    g599(.A(new_n635), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n553), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n727), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n727), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n656), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(G85gat), .B1(new_n808), .B2(new_n458), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n801), .A2(new_n553), .A3(new_n769), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n711), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n463), .A2(new_n425), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  NAND3_X1  g612(.A1(new_n711), .A2(new_n459), .A3(new_n810), .ZN(new_n814));
  INV_X1    g613(.A(new_n557), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n459), .A2(new_n564), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n816), .B(new_n820), .C1(new_n807), .C2(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT120), .B(G99gat), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n399), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n811), .A2(new_n674), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n823), .ZN(G1338gat));
  NAND3_X1  g626(.A1(new_n811), .A2(G106gat), .A3(new_n283), .ZN(new_n828));
  INV_X1    g627(.A(G106gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n807), .B2(new_n443), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1339gat));
  NAND4_X1  g634(.A1(new_n553), .A2(new_n608), .A3(new_n769), .A4(new_n635), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n621), .A2(new_n618), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n617), .A2(new_n619), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n627), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n656), .A2(new_n632), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n646), .B(new_n642), .C1(new_n645), .C2(KEYINPUT10), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n636), .C1(new_n641), .C2(new_n643), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n653), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n841), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n644), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n653), .A4(new_n845), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n655), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n840), .B1(new_n850), .B2(new_n635), .ZN(new_n851));
  INV_X1    g650(.A(new_n850), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n839), .A2(new_n632), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n604), .B2(new_n607), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n851), .A2(new_n608), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n836), .B1(new_n855), .B2(new_n553), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(new_n443), .A3(new_n399), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n463), .A2(new_n459), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n635), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n856), .A2(new_n767), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n717), .A2(new_n362), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n635), .A2(G113gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  OAI21_X1  g666(.A(G120gat), .B1(new_n860), .B2(new_n769), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n769), .A2(G120gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n865), .B2(new_n869), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n859), .A2(G127gat), .A3(new_n553), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT121), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT121), .ZN(new_n873));
  INV_X1    g672(.A(new_n865), .ZN(new_n874));
  AOI21_X1  g673(.A(G127gat), .B1(new_n874), .B2(new_n553), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(G1342gat));
  OR3_X1    g675(.A1(new_n865), .A2(G134gat), .A3(new_n608), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n860), .B2(new_n608), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n856), .A2(new_n882), .A3(new_n283), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n856), .B2(new_n283), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n478), .A2(new_n858), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G141gat), .B1(new_n887), .B2(new_n635), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n674), .A2(new_n443), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n862), .A2(new_n362), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n236), .A3(new_n801), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n226), .A3(new_n656), .ZN(new_n894));
  INV_X1    g693(.A(new_n887), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT59), .B(new_n226), .C1(new_n895), .C2(new_n656), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n443), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n883), .B2(new_n884), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n856), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n443), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n900), .A2(new_n656), .A3(new_n886), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n894), .B1(new_n896), .B2(new_n904), .ZN(G1345gat));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n553), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n907));
  AOI21_X1  g706(.A(G155gat), .B1(new_n906), .B2(KEYINPUT123), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n553), .A2(G155gat), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n907), .A2(new_n908), .B1(new_n895), .B2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n887), .B2(new_n608), .ZN(new_n911));
  INV_X1    g710(.A(G162gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n912), .A3(new_n609), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1347gat));
  AND3_X1   g713(.A1(new_n856), .A2(new_n463), .A3(new_n459), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(new_n717), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n296), .A3(new_n801), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n767), .A2(new_n362), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n857), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n635), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT124), .Z(G1348gat));
  AOI21_X1  g721(.A(G176gat), .B1(new_n916), .B2(new_n656), .ZN(new_n923));
  INV_X1    g722(.A(new_n919), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n769), .A2(new_n304), .A3(new_n305), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G1349gat));
  OAI211_X1 g725(.A(new_n916), .B(new_n553), .C1(new_n317), .C2(new_n316), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n919), .B2(new_n554), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n919), .B2(new_n608), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n310), .A3(new_n609), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n889), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n935), .A2(G197gat), .A3(new_n635), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n856), .A2(new_n283), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT57), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n856), .A2(new_n882), .A3(new_n283), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n898), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n940), .B2(new_n901), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n900), .A2(new_n942), .A3(new_n902), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n673), .A2(new_n918), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n941), .A2(new_n801), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT126), .ZN(new_n946));
  OAI21_X1  g745(.A(G197gat), .B1(new_n945), .B2(KEYINPUT126), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n936), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n949), .B2(new_n769), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n935), .A2(G204gat), .A3(new_n769), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  OR3_X1    g752(.A1(new_n935), .A2(G211gat), .A3(new_n554), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n944), .A2(new_n553), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n900), .A2(new_n902), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(KEYINPUT127), .B(new_n954), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1354gat));
  INV_X1    g762(.A(G218gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n949), .A2(new_n964), .A3(new_n608), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n915), .A2(new_n609), .A3(new_n889), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(G1355gat));
endmodule


