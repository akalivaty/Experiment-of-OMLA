

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778;

  NOR2_X1 U369 ( .A1(G953), .A2(G237), .ZN(n538) );
  NOR2_X1 U370 ( .A1(n736), .A2(n735), .ZN(n347) );
  NOR2_X1 U371 ( .A1(n719), .A2(n718), .ZN(n642) );
  XNOR2_X2 U372 ( .A(n430), .B(n551), .ZN(n611) );
  NOR2_X2 U373 ( .A1(n508), .A2(n456), .ZN(n441) );
  XNOR2_X2 U374 ( .A(n412), .B(KEYINPUT46), .ZN(n508) );
  NOR2_X1 U375 ( .A1(n718), .A2(n411), .ZN(n646) );
  XNOR2_X1 U376 ( .A(n411), .B(n524), .ZN(n719) );
  XNOR2_X2 U377 ( .A(n592), .B(KEYINPUT80), .ZN(n683) );
  XNOR2_X2 U378 ( .A(n644), .B(n495), .ZN(n640) );
  BUF_X2 U379 ( .A(n738), .Z(n748) );
  NOR2_X1 U380 ( .A1(n410), .A2(n675), .ZN(n408) );
  XNOR2_X1 U381 ( .A(n416), .B(n415), .ZN(n434) );
  XNOR2_X1 U382 ( .A(n516), .B(n506), .ZN(n375) );
  AND2_X1 U383 ( .A1(n368), .A2(n367), .ZN(n366) );
  NOR2_X1 U384 ( .A1(n683), .A2(n596), .ZN(n597) );
  XNOR2_X1 U385 ( .A(n375), .B(n388), .ZN(n703) );
  AND2_X1 U386 ( .A1(n429), .A2(n612), .ZN(n684) );
  INV_X1 U387 ( .A(n611), .ZN(n429) );
  NOR2_X1 U388 ( .A1(n663), .A2(G902), .ZN(n430) );
  INV_X1 U389 ( .A(KEYINPUT85), .ZN(n654) );
  XNOR2_X1 U390 ( .A(n361), .B(KEYINPUT119), .ZN(n360) );
  AND2_X2 U391 ( .A1(n369), .A2(n366), .ZN(n365) );
  NAND2_X1 U392 ( .A1(n766), .A2(n370), .ZN(n368) );
  OR2_X1 U393 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U394 ( .A(n406), .B(n405), .ZN(n648) );
  NOR2_X1 U395 ( .A1(n737), .A2(n347), .ZN(n372) );
  AND2_X1 U396 ( .A1(n414), .A2(n409), .ZN(n675) );
  AND2_X1 U397 ( .A1(n697), .A2(n394), .ZN(n420) );
  AND2_X1 U398 ( .A1(n404), .A2(n647), .ZN(n410) );
  NAND2_X1 U399 ( .A1(n620), .A2(KEYINPUT86), .ZN(n454) );
  NAND2_X1 U400 ( .A1(n417), .A2(n436), .ZN(n416) );
  XNOR2_X1 U401 ( .A(n597), .B(KEYINPUT73), .ZN(n419) );
  AND2_X1 U402 ( .A1(n609), .A2(n598), .ZN(n394) );
  XNOR2_X1 U403 ( .A(n481), .B(n389), .ZN(n417) );
  AND2_X1 U404 ( .A1(n402), .A2(n469), .ZN(n643) );
  AND2_X1 U405 ( .A1(n622), .A2(n688), .ZN(n618) );
  AND2_X1 U406 ( .A1(n355), .A2(n353), .ZN(n352) );
  NOR2_X1 U407 ( .A1(n437), .A2(n705), .ZN(n614) );
  XNOR2_X1 U408 ( .A(n349), .B(KEYINPUT110), .ZN(n437) );
  NAND2_X1 U409 ( .A1(n703), .A2(n702), .ZN(n349) );
  NOR2_X1 U410 ( .A1(n385), .A2(n354), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n584), .B(n583), .ZN(n589) );
  OR2_X1 U412 ( .A1(n705), .A2(n629), .ZN(n385) );
  AND2_X1 U413 ( .A1(n627), .A2(n470), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n557), .B(n556), .ZN(n612) );
  NOR2_X1 U415 ( .A1(G902), .A2(n657), .ZN(n523) );
  XNOR2_X1 U416 ( .A(n514), .B(n513), .ZN(n515) );
  BUF_X1 U417 ( .A(n519), .Z(n477) );
  NOR2_X1 U418 ( .A1(n371), .A2(n654), .ZN(n370) );
  XNOR2_X1 U419 ( .A(n554), .B(n504), .ZN(n519) );
  XNOR2_X1 U420 ( .A(n546), .B(G134), .ZN(n464) );
  XNOR2_X1 U421 ( .A(n486), .B(G104), .ZN(n545) );
  XNOR2_X1 U422 ( .A(n487), .B(G110), .ZN(n567) );
  XNOR2_X1 U423 ( .A(n505), .B(G143), .ZN(n554) );
  INV_X1 U424 ( .A(n655), .ZN(n371) );
  INV_X2 U425 ( .A(KEYINPUT3), .ZN(n484) );
  XNOR2_X1 U426 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n509) );
  INV_X2 U427 ( .A(KEYINPUT67), .ZN(n480) );
  NAND2_X1 U428 ( .A1(n348), .A2(n413), .ZN(n412) );
  XNOR2_X2 U429 ( .A(n483), .B(KEYINPUT42), .ZN(n348) );
  XNOR2_X1 U430 ( .A(n348), .B(G137), .ZN(G39) );
  INV_X1 U431 ( .A(n377), .ZN(n364) );
  NOR2_X2 U432 ( .A1(n377), .A2(n766), .ZN(n374) );
  NAND2_X1 U433 ( .A1(n377), .A2(n370), .ZN(n369) );
  XNOR2_X2 U434 ( .A(n498), .B(n497), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n403), .A2(n627), .ZN(n628) );
  NAND2_X1 U436 ( .A1(n352), .A2(n350), .ZN(n481) );
  NAND2_X1 U437 ( .A1(n403), .A2(n351), .ZN(n350) );
  NOR2_X1 U438 ( .A1(n627), .A2(n470), .ZN(n354) );
  NAND2_X1 U439 ( .A1(n356), .A2(KEYINPUT0), .ZN(n355) );
  INV_X1 U440 ( .A(n403), .ZN(n356) );
  XNOR2_X2 U441 ( .A(n588), .B(KEYINPUT19), .ZN(n403) );
  XNOR2_X1 U442 ( .A(n358), .B(n357), .ZN(G75) );
  INV_X1 U443 ( .A(KEYINPUT53), .ZN(n357) );
  NAND2_X1 U444 ( .A1(n360), .A2(n359), .ZN(n358) );
  INV_X1 U445 ( .A(G953), .ZN(n359) );
  NAND2_X1 U446 ( .A1(n373), .A2(n372), .ZN(n361) );
  NAND2_X1 U447 ( .A1(n365), .A2(n362), .ZN(n435) );
  NAND2_X1 U448 ( .A1(n364), .A2(n363), .ZN(n362) );
  NOR2_X1 U449 ( .A1(n766), .A2(n655), .ZN(n363) );
  NAND2_X1 U450 ( .A1(n371), .A2(n654), .ZN(n367) );
  NAND2_X2 U451 ( .A1(n482), .A2(n700), .ZN(n766) );
  XNOR2_X1 U452 ( .A(n734), .B(n733), .ZN(n373) );
  XNOR2_X1 U453 ( .A(n516), .B(n506), .ZN(n610) );
  XNOR2_X1 U454 ( .A(n484), .B(G116), .ZN(n376) );
  XNOR2_X1 U455 ( .A(n471), .B(n525), .ZN(n378) );
  INV_X1 U456 ( .A(KEYINPUT4), .ZN(n504) );
  OR2_X1 U457 ( .A1(G237), .A2(G902), .ZN(n558) );
  NOR2_X1 U458 ( .A1(n379), .A2(n440), .ZN(n439) );
  AND2_X1 U459 ( .A1(n619), .A2(n456), .ZN(n379) );
  NAND2_X1 U460 ( .A1(n455), .A2(n496), .ZN(n440) );
  NAND2_X1 U461 ( .A1(n452), .A2(n496), .ZN(n451) );
  INV_X1 U462 ( .A(KEYINPUT8), .ZN(n489) );
  INV_X1 U463 ( .A(KEYINPUT69), .ZN(n583) );
  INV_X1 U464 ( .A(KEYINPUT6), .ZN(n495) );
  INV_X1 U465 ( .A(n604), .ZN(n467) );
  OR2_X2 U466 ( .A1(n711), .A2(n629), .ZN(n718) );
  INV_X1 U467 ( .A(KEYINPUT0), .ZN(n470) );
  XNOR2_X1 U468 ( .A(n485), .B(n567), .ZN(n473) );
  XNOR2_X1 U469 ( .A(n509), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U470 ( .A(KEYINPUT9), .B(KEYINPUT103), .ZN(n553) );
  XNOR2_X1 U471 ( .A(n552), .B(n424), .ZN(n423) );
  XNOR2_X1 U472 ( .A(G134), .B(G116), .ZN(n552) );
  XNOR2_X1 U473 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n424) );
  XNOR2_X1 U474 ( .A(n463), .B(n462), .ZN(n461) );
  XNOR2_X1 U475 ( .A(n384), .B(n518), .ZN(n462) );
  XNOR2_X1 U476 ( .A(n517), .B(n572), .ZN(n463) );
  XNOR2_X1 U477 ( .A(n555), .B(G478), .ZN(n556) );
  NOR2_X1 U478 ( .A1(G902), .A2(n746), .ZN(n557) );
  BUF_X1 U479 ( .A(n711), .Z(n433) );
  XOR2_X1 U480 ( .A(KEYINPUT92), .B(n661), .Z(n744) );
  INV_X1 U481 ( .A(KEYINPUT88), .ZN(n405) );
  INV_X1 U482 ( .A(n515), .ZN(n390) );
  INV_X2 U483 ( .A(G128), .ZN(n505) );
  INV_X1 U484 ( .A(G113), .ZN(n486) );
  XNOR2_X1 U485 ( .A(G143), .B(G122), .ZN(n541) );
  XOR2_X1 U486 ( .A(KEYINPUT11), .B(G140), .Z(n542) );
  XOR2_X1 U487 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n540) );
  XOR2_X1 U488 ( .A(G137), .B(G140), .Z(n572) );
  XNOR2_X1 U489 ( .A(G902), .B(KEYINPUT15), .ZN(n655) );
  XOR2_X1 U490 ( .A(KEYINPUT66), .B(G101), .Z(n520) );
  XOR2_X1 U491 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n511) );
  NAND2_X1 U492 ( .A1(G234), .A2(G237), .ZN(n575) );
  XNOR2_X1 U493 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U494 ( .A(G137), .B(G119), .ZN(n526) );
  NAND2_X1 U495 ( .A1(n439), .A2(n438), .ZN(n449) );
  INV_X1 U496 ( .A(KEYINPUT45), .ZN(n497) );
  INV_X1 U497 ( .A(KEYINPUT23), .ZN(n564) );
  INV_X1 U498 ( .A(G119), .ZN(n487) );
  INV_X1 U499 ( .A(KEYINPUT33), .ZN(n493) );
  XNOR2_X1 U500 ( .A(n684), .B(n428), .ZN(n621) );
  INV_X1 U501 ( .A(KEYINPUT105), .ZN(n428) );
  NAND2_X1 U502 ( .A1(n380), .A2(n466), .ZN(n617) );
  XNOR2_X1 U503 ( .A(n425), .B(n421), .ZN(n746) );
  XNOR2_X1 U504 ( .A(n423), .B(n422), .ZN(n421) );
  XNOR2_X1 U505 ( .A(n553), .B(KEYINPUT101), .ZN(n422) );
  XNOR2_X1 U506 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n600) );
  INV_X1 U507 ( .A(n723), .ZN(n469) );
  INV_X1 U508 ( .A(n612), .ZN(n593) );
  NOR2_X1 U509 ( .A1(n640), .A2(n433), .ZN(n409) );
  XNOR2_X1 U510 ( .A(n660), .B(n507), .ZN(n662) );
  INV_X1 U511 ( .A(KEYINPUT56), .ZN(n500) );
  XOR2_X1 U512 ( .A(KEYINPUT30), .B(n603), .Z(n380) );
  XNOR2_X1 U513 ( .A(n641), .B(KEYINPUT77), .ZN(n381) );
  AND2_X1 U514 ( .A1(n636), .A2(n635), .ZN(n382) );
  NOR2_X1 U515 ( .A1(n619), .A2(n454), .ZN(n383) );
  BUF_X1 U516 ( .A(n719), .Z(n436) );
  XOR2_X1 U517 ( .A(G104), .B(G110), .Z(n384) );
  AND2_X1 U518 ( .A1(n453), .A2(n456), .ZN(n386) );
  XNOR2_X1 U519 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n387) );
  XNOR2_X1 U520 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n388) );
  XOR2_X1 U521 ( .A(KEYINPUT22), .B(KEYINPUT64), .Z(n389) );
  INV_X1 U522 ( .A(KEYINPUT48), .ZN(n456) );
  INV_X1 U523 ( .A(KEYINPUT86), .ZN(n496) );
  INV_X1 U524 ( .A(KEYINPUT2), .ZN(n733) );
  XNOR2_X1 U525 ( .A(n397), .B(n390), .ZN(n742) );
  XNOR2_X2 U526 ( .A(n478), .B(n477), .ZN(n397) );
  INV_X1 U527 ( .A(n545), .ZN(n475) );
  NAND2_X1 U528 ( .A1(n378), .A2(n475), .ZN(n392) );
  NAND2_X1 U529 ( .A1(n391), .A2(n545), .ZN(n393) );
  NAND2_X1 U530 ( .A1(n393), .A2(n392), .ZN(n474) );
  INV_X1 U531 ( .A(n476), .ZN(n391) );
  XNOR2_X1 U532 ( .A(n471), .B(n525), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U534 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U535 ( .A(n505), .B(G143), .ZN(n395) );
  NAND2_X1 U536 ( .A1(n434), .A2(n630), .ZN(n396) );
  NAND2_X1 U537 ( .A1(n434), .A2(n630), .ZN(n632) );
  XNOR2_X1 U538 ( .A(n637), .B(KEYINPUT78), .ZN(n638) );
  NOR2_X1 U539 ( .A1(n671), .A2(G902), .ZN(n537) );
  INV_X1 U540 ( .A(n397), .ZN(n398) );
  NAND2_X1 U541 ( .A1(n693), .A2(n678), .ZN(n404) );
  XNOR2_X1 U542 ( .A(n396), .B(n631), .ZN(n399) );
  BUF_X1 U543 ( .A(n478), .Z(n400) );
  XNOR2_X1 U544 ( .A(n632), .B(n631), .ZN(n479) );
  XOR2_X1 U545 ( .A(n671), .B(KEYINPUT62), .Z(n673) );
  AND2_X1 U546 ( .A1(n445), .A2(n444), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n398), .B(n515), .ZN(n401) );
  NAND2_X1 U548 ( .A1(n508), .A2(n456), .ZN(n455) );
  AND2_X1 U549 ( .A1(n646), .A2(n467), .ZN(n466) );
  OR2_X2 U550 ( .A1(n750), .A2(G902), .ZN(n492) );
  NAND2_X1 U551 ( .A1(n776), .A2(KEYINPUT44), .ZN(n407) );
  NAND2_X1 U552 ( .A1(n431), .A2(n744), .ZN(n674) );
  XNOR2_X1 U553 ( .A(n672), .B(n673), .ZN(n431) );
  NAND2_X1 U554 ( .A1(n502), .A2(n744), .ZN(n501) );
  XNOR2_X1 U555 ( .A(n503), .B(n743), .ZN(n502) );
  XNOR2_X2 U556 ( .A(n628), .B(n470), .ZN(n402) );
  NAND2_X1 U557 ( .A1(n615), .A2(n403), .ZN(n592) );
  NAND2_X1 U558 ( .A1(n645), .A2(n646), .ZN(n678) );
  XNOR2_X2 U559 ( .A(n643), .B(KEYINPUT31), .ZN(n693) );
  NOR2_X1 U560 ( .A1(n591), .A2(n411), .ZN(n615) );
  XNOR2_X2 U561 ( .A(n523), .B(G469), .ZN(n411) );
  XNOR2_X2 U562 ( .A(n492), .B(n574), .ZN(n711) );
  INV_X1 U563 ( .A(n777), .ZN(n413) );
  INV_X1 U564 ( .A(n416), .ZN(n414) );
  INV_X1 U565 ( .A(KEYINPUT108), .ZN(n415) );
  NAND2_X1 U566 ( .A1(n417), .A2(n382), .ZN(n637) );
  XNOR2_X2 U567 ( .A(n418), .B(KEYINPUT68), .ZN(n619) );
  NAND2_X1 U568 ( .A1(n420), .A2(n419), .ZN(n418) );
  XNOR2_X1 U569 ( .A(n427), .B(n426), .ZN(n425) );
  XNOR2_X1 U570 ( .A(n395), .B(n471), .ZN(n426) );
  XNOR2_X2 U571 ( .A(n472), .B(G122), .ZN(n471) );
  NAND2_X1 U572 ( .A1(n563), .A2(G217), .ZN(n427) );
  XNOR2_X2 U573 ( .A(n490), .B(n489), .ZN(n563) );
  NAND2_X1 U574 ( .A1(n468), .A2(n402), .ZN(n460) );
  AND2_X1 U575 ( .A1(n402), .A2(n716), .ZN(n645) );
  NAND2_X2 U576 ( .A1(n642), .A2(n640), .ZN(n494) );
  INV_X2 U577 ( .A(G107), .ZN(n472) );
  XNOR2_X1 U578 ( .A(n432), .B(n590), .ZN(n591) );
  NOR2_X1 U579 ( .A1(n589), .A2(n716), .ZN(n432) );
  XNOR2_X1 U580 ( .A(n374), .B(n733), .ZN(n656) );
  AND2_X2 U581 ( .A1(n435), .A2(n656), .ZN(n738) );
  NOR2_X1 U582 ( .A1(n706), .A2(n437), .ZN(n707) );
  INV_X1 U583 ( .A(n619), .ZN(n442) );
  NAND2_X1 U584 ( .A1(n441), .A2(n442), .ZN(n438) );
  NAND2_X1 U585 ( .A1(n383), .A2(n441), .ZN(n444) );
  AND2_X1 U586 ( .A1(n619), .A2(n443), .ZN(n446) );
  NOR2_X1 U587 ( .A1(n454), .A2(KEYINPUT48), .ZN(n443) );
  NAND2_X1 U588 ( .A1(n386), .A2(n508), .ZN(n448) );
  NOR2_X1 U589 ( .A1(n447), .A2(n446), .ZN(n445) );
  NAND2_X1 U590 ( .A1(n448), .A2(n451), .ZN(n447) );
  NAND2_X1 U591 ( .A1(n450), .A2(n449), .ZN(n482) );
  INV_X1 U592 ( .A(n620), .ZN(n452) );
  INV_X1 U593 ( .A(n454), .ZN(n453) );
  XNOR2_X2 U594 ( .A(n457), .B(n387), .ZN(n776) );
  NAND2_X1 U595 ( .A1(n458), .A2(n381), .ZN(n457) );
  XNOR2_X1 U596 ( .A(n460), .B(n459), .ZN(n458) );
  INV_X1 U597 ( .A(KEYINPUT34), .ZN(n459) );
  XNOR2_X1 U598 ( .A(n533), .B(n461), .ZN(n657) );
  XNOR2_X2 U599 ( .A(n765), .B(n522), .ZN(n533) );
  XNOR2_X2 U600 ( .A(n519), .B(n464), .ZN(n765) );
  XNOR2_X1 U601 ( .A(n465), .B(n491), .ZN(n622) );
  NOR2_X2 U602 ( .A1(n617), .A2(n616), .ZN(n465) );
  INV_X1 U603 ( .A(n735), .ZN(n468) );
  XNOR2_X2 U604 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n400), .B(G101), .ZN(n759) );
  NAND2_X1 U606 ( .A1(n479), .A2(n775), .ZN(n652) );
  XNOR2_X1 U607 ( .A(n399), .B(G110), .ZN(G12) );
  XNOR2_X2 U608 ( .A(n480), .B(G131), .ZN(n546) );
  XOR2_X2 U609 ( .A(KEYINPUT106), .B(n595), .Z(n706) );
  XOR2_X2 U610 ( .A(G146), .B(G125), .Z(n547) );
  XNOR2_X1 U611 ( .A(n573), .B(n764), .ZN(n750) );
  INV_X1 U612 ( .A(n703), .ZN(n616) );
  NAND2_X1 U613 ( .A1(n710), .A2(n615), .ZN(n483) );
  XNOR2_X2 U614 ( .A(n484), .B(G116), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n566), .B(n488), .ZN(n569) );
  NAND2_X1 U616 ( .A1(n563), .A2(G221), .ZN(n488) );
  NAND2_X1 U617 ( .A1(n758), .A2(G234), .ZN(n490) );
  INV_X1 U618 ( .A(KEYINPUT39), .ZN(n491) );
  XNOR2_X2 U619 ( .A(n494), .B(n493), .ZN(n735) );
  NAND2_X1 U620 ( .A1(n499), .A2(n653), .ZN(n498) );
  XNOR2_X1 U621 ( .A(n650), .B(KEYINPUT87), .ZN(n499) );
  XNOR2_X1 U622 ( .A(n501), .B(n500), .ZN(G51) );
  NAND2_X1 U623 ( .A1(n738), .A2(G210), .ZN(n503) );
  AND2_X1 U624 ( .A1(G210), .A2(n558), .ZN(n506) );
  XOR2_X1 U625 ( .A(n659), .B(n658), .Z(n507) );
  OR2_X1 U626 ( .A1(n706), .A2(KEYINPUT47), .ZN(n596) );
  XNOR2_X1 U627 ( .A(n521), .B(G146), .ZN(n522) );
  INV_X1 U628 ( .A(KEYINPUT104), .ZN(n555) );
  XNOR2_X1 U629 ( .A(n535), .B(G472), .ZN(n536) );
  XNOR2_X1 U630 ( .A(KEYINPUT13), .B(G475), .ZN(n551) );
  XNOR2_X1 U631 ( .A(n601), .B(n600), .ZN(n602) );
  BUF_X1 U632 ( .A(n375), .Z(n606) );
  INV_X1 U633 ( .A(KEYINPUT60), .ZN(n669) );
  NOR2_X1 U634 ( .A1(n662), .A2(n752), .ZN(G54) );
  INV_X2 U635 ( .A(G953), .ZN(n758) );
  NAND2_X1 U636 ( .A1(G224), .A2(n758), .ZN(n510) );
  XNOR2_X1 U637 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U638 ( .A(n512), .B(KEYINPUT90), .Z(n514) );
  XNOR2_X1 U639 ( .A(n520), .B(n547), .ZN(n513) );
  NAND2_X1 U640 ( .A1(n742), .A2(n655), .ZN(n516) );
  XOR2_X1 U641 ( .A(KEYINPUT94), .B(G107), .Z(n517) );
  NAND2_X1 U642 ( .A1(G227), .A2(n758), .ZN(n518) );
  INV_X1 U643 ( .A(n520), .ZN(n521) );
  XOR2_X1 U644 ( .A(KEYINPUT65), .B(KEYINPUT1), .Z(n524) );
  XNOR2_X1 U645 ( .A(n526), .B(n376), .ZN(n530) );
  XOR2_X1 U646 ( .A(G113), .B(KEYINPUT98), .Z(n528) );
  XNOR2_X1 U647 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U648 ( .A(n530), .B(n529), .Z(n532) );
  NAND2_X1 U649 ( .A1(n538), .A2(G210), .ZN(n531) );
  XNOR2_X1 U650 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U651 ( .A(n534), .B(n533), .ZN(n671) );
  XNOR2_X1 U652 ( .A(KEYINPUT99), .B(KEYINPUT70), .ZN(n535) );
  XNOR2_X2 U653 ( .A(n537), .B(n536), .ZN(n644) );
  INV_X1 U654 ( .A(n640), .ZN(n639) );
  NAND2_X1 U655 ( .A1(G214), .A2(n538), .ZN(n539) );
  XNOR2_X1 U656 ( .A(n540), .B(n539), .ZN(n544) );
  XNOR2_X1 U657 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U658 ( .A(n544), .B(n543), .Z(n550) );
  XNOR2_X1 U659 ( .A(n546), .B(n545), .ZN(n548) );
  XNOR2_X1 U660 ( .A(n547), .B(KEYINPUT10), .ZN(n570) );
  XNOR2_X1 U661 ( .A(n548), .B(n570), .ZN(n549) );
  XNOR2_X1 U662 ( .A(n550), .B(n549), .ZN(n663) );
  NAND2_X1 U663 ( .A1(n611), .A2(n593), .ZN(n691) );
  INV_X1 U664 ( .A(n691), .ZN(n688) );
  NAND2_X1 U665 ( .A1(G214), .A2(n558), .ZN(n702) );
  NAND2_X1 U666 ( .A1(n688), .A2(n702), .ZN(n559) );
  OR2_X1 U667 ( .A1(n639), .A2(n559), .ZN(n585) );
  XOR2_X1 U668 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n562) );
  NAND2_X1 U669 ( .A1(n655), .A2(G234), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n560), .B(KEYINPUT20), .ZN(n580) );
  NAND2_X1 U671 ( .A1(n580), .A2(G217), .ZN(n561) );
  XNOR2_X1 U672 ( .A(n562), .B(n561), .ZN(n574) );
  XOR2_X1 U673 ( .A(G128), .B(KEYINPUT84), .Z(n565) );
  XNOR2_X1 U674 ( .A(n567), .B(KEYINPUT24), .ZN(n568) );
  XNOR2_X1 U675 ( .A(n569), .B(n568), .ZN(n573) );
  INV_X1 U676 ( .A(n570), .ZN(n571) );
  XNOR2_X1 U677 ( .A(n572), .B(n571), .ZN(n764) );
  XNOR2_X1 U678 ( .A(n575), .B(KEYINPUT14), .ZN(n576) );
  XNOR2_X1 U679 ( .A(KEYINPUT74), .B(n576), .ZN(n577) );
  NAND2_X1 U680 ( .A1(G952), .A2(n577), .ZN(n732) );
  NOR2_X1 U681 ( .A1(G953), .A2(n732), .ZN(n625) );
  AND2_X1 U682 ( .A1(n577), .A2(G953), .ZN(n578) );
  NAND2_X1 U683 ( .A1(G902), .A2(n578), .ZN(n623) );
  NOR2_X1 U684 ( .A1(G900), .A2(n623), .ZN(n579) );
  NOR2_X1 U685 ( .A1(n625), .A2(n579), .ZN(n604) );
  NAND2_X1 U686 ( .A1(G221), .A2(n580), .ZN(n581) );
  XNOR2_X1 U687 ( .A(KEYINPUT21), .B(n581), .ZN(n712) );
  NOR2_X1 U688 ( .A1(n604), .A2(n712), .ZN(n582) );
  NAND2_X1 U689 ( .A1(n711), .A2(n582), .ZN(n584) );
  NOR2_X1 U690 ( .A1(n585), .A2(n589), .ZN(n599) );
  AND2_X1 U691 ( .A1(n436), .A2(n599), .ZN(n586) );
  XNOR2_X1 U692 ( .A(n586), .B(KEYINPUT43), .ZN(n587) );
  NOR2_X1 U693 ( .A1(n606), .A2(n587), .ZN(n701) );
  INV_X1 U694 ( .A(n701), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n610), .A2(n702), .ZN(n588) );
  INV_X1 U696 ( .A(KEYINPUT28), .ZN(n590) );
  INV_X1 U697 ( .A(n644), .ZN(n716) );
  INV_X1 U698 ( .A(n621), .ZN(n594) );
  NAND2_X1 U699 ( .A1(n691), .A2(n594), .ZN(n595) );
  NAND2_X1 U700 ( .A1(n683), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U701 ( .A1(n599), .A2(n606), .ZN(n601) );
  XNOR2_X1 U702 ( .A(n719), .B(KEYINPUT91), .ZN(n633) );
  NAND2_X1 U703 ( .A1(n602), .A2(n633), .ZN(n697) );
  NAND2_X1 U704 ( .A1(KEYINPUT47), .A2(n706), .ZN(n607) );
  XNOR2_X1 U705 ( .A(KEYINPUT96), .B(n712), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n644), .A2(n702), .ZN(n603) );
  NAND2_X1 U707 ( .A1(n611), .A2(n612), .ZN(n641) );
  NOR2_X1 U708 ( .A1(n617), .A2(n641), .ZN(n605) );
  NAND2_X1 U709 ( .A1(n606), .A2(n605), .ZN(n687) );
  NAND2_X1 U710 ( .A1(n607), .A2(n687), .ZN(n608) );
  XNOR2_X1 U711 ( .A(n608), .B(KEYINPUT81), .ZN(n609) );
  OR2_X1 U712 ( .A1(n612), .A2(n611), .ZN(n705) );
  XNOR2_X1 U713 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n613) );
  XNOR2_X1 U714 ( .A(n614), .B(n613), .ZN(n710) );
  XNOR2_X1 U715 ( .A(KEYINPUT40), .B(n618), .ZN(n777) );
  NAND2_X1 U716 ( .A1(n622), .A2(n621), .ZN(n700) );
  NOR2_X1 U717 ( .A1(G898), .A2(n623), .ZN(n624) );
  NOR2_X1 U718 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U719 ( .A(KEYINPUT93), .B(n626), .ZN(n627) );
  AND2_X1 U720 ( .A1(n716), .A2(n433), .ZN(n630) );
  INV_X1 U721 ( .A(KEYINPUT109), .ZN(n631) );
  XNOR2_X1 U722 ( .A(n640), .B(KEYINPUT79), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n633), .A2(n433), .ZN(n634) );
  XNOR2_X1 U724 ( .A(KEYINPUT107), .B(n634), .ZN(n635) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U726 ( .A1(n652), .A2(KEYINPUT44), .ZN(n649) );
  INV_X1 U727 ( .A(n706), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n642), .A2(n644), .ZN(n723) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  OR2_X1 U730 ( .A1(n776), .A2(KEYINPUT44), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n748), .A2(G469), .ZN(n660) );
  XOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n659) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT121), .ZN(n658) );
  NOR2_X1 U734 ( .A1(G952), .A2(n758), .ZN(n661) );
  INV_X1 U735 ( .A(n744), .ZN(n752) );
  NAND2_X1 U736 ( .A1(n738), .A2(G475), .ZN(n667) );
  XOR2_X1 U737 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n665) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT122), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n668), .A2(n744), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n738), .A2(G472), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U745 ( .A(G101), .B(n675), .Z(G3) );
  NOR2_X1 U746 ( .A1(n691), .A2(n678), .ZN(n676) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(n676), .Z(n677) );
  XNOR2_X1 U748 ( .A(G104), .B(n677), .ZN(G6) );
  INV_X1 U749 ( .A(n684), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n678), .A2(n694), .ZN(n682) );
  XOR2_X1 U751 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n680) );
  XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT27), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n682), .B(n681), .ZN(G9) );
  XOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .Z(n686) );
  INV_X1 U756 ( .A(n683), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n684), .A2(n689), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(G30) );
  XNOR2_X1 U759 ( .A(G143), .B(n687), .ZN(G45) );
  NAND2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n690), .B(G146), .ZN(G48) );
  NOR2_X1 U762 ( .A1(n691), .A2(n693), .ZN(n692) );
  XOR2_X1 U763 ( .A(G113), .B(n692), .Z(G15) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U765 ( .A(KEYINPUT114), .B(n695), .Z(n696) );
  XNOR2_X1 U766 ( .A(G116), .B(n696), .ZN(G18) );
  XNOR2_X1 U767 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n698) );
  XNOR2_X1 U768 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U769 ( .A(G125), .B(n699), .ZN(G27) );
  XNOR2_X1 U770 ( .A(G134), .B(n700), .ZN(G36) );
  XOR2_X1 U771 ( .A(G140), .B(n701), .Z(G42) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U775 ( .A1(n709), .A2(n735), .ZN(n728) );
  INV_X1 U776 ( .A(n710), .ZN(n736) );
  XOR2_X1 U777 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n714) );
  NAND2_X1 U778 ( .A1(n712), .A2(n433), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U781 ( .A(n717), .B(KEYINPUT117), .ZN(n722) );
  NAND2_X1 U782 ( .A1(n436), .A2(n718), .ZN(n720) );
  XNOR2_X1 U783 ( .A(KEYINPUT50), .B(n720), .ZN(n721) );
  NAND2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U785 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U786 ( .A(KEYINPUT51), .B(n725), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n736), .A2(n726), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U789 ( .A(n729), .B(KEYINPUT52), .ZN(n730) );
  XNOR2_X1 U790 ( .A(KEYINPUT118), .B(n730), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n374), .A2(KEYINPUT83), .ZN(n734) );
  XOR2_X1 U793 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n740) );
  XNOR2_X1 U794 ( .A(KEYINPUT82), .B(KEYINPUT55), .ZN(n739) );
  XNOR2_X1 U795 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n401), .B(n741), .ZN(n743) );
  NAND2_X1 U797 ( .A1(G478), .A2(n748), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n745), .B(n746), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n747), .A2(n752), .ZN(G63) );
  NAND2_X1 U800 ( .A1(G217), .A2(n748), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n749), .B(n750), .ZN(n751) );
  NOR2_X1 U802 ( .A1(n751), .A2(n752), .ZN(G66) );
  INV_X1 U803 ( .A(G898), .ZN(n755) );
  NAND2_X1 U804 ( .A1(G953), .A2(G224), .ZN(n753) );
  XOR2_X1 U805 ( .A(KEYINPUT61), .B(n753), .Z(n754) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n757) );
  NOR2_X1 U807 ( .A1(G953), .A2(n377), .ZN(n756) );
  NOR2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n763) );
  NOR2_X1 U809 ( .A1(G898), .A2(n758), .ZN(n760) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U811 ( .A(KEYINPUT124), .B(n761), .Z(n762) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(G69) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(n769) );
  XOR2_X1 U814 ( .A(n766), .B(n769), .Z(n767) );
  NOR2_X1 U815 ( .A1(G953), .A2(n767), .ZN(n768) );
  XNOR2_X1 U816 ( .A(KEYINPUT125), .B(n768), .ZN(n774) );
  XNOR2_X1 U817 ( .A(G227), .B(n769), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G953), .ZN(n772) );
  XNOR2_X1 U820 ( .A(KEYINPUT126), .B(n772), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(G72) );
  XNOR2_X1 U822 ( .A(G119), .B(n775), .ZN(G21) );
  XOR2_X1 U823 ( .A(n776), .B(G122), .Z(G24) );
  XNOR2_X1 U824 ( .A(G131), .B(KEYINPUT127), .ZN(n778) );
  XNOR2_X1 U825 ( .A(n778), .B(n777), .ZN(G33) );
endmodule

