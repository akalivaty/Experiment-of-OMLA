//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n478), .A2(new_n482), .A3(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n474), .B2(new_n475), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(new_n490), .C1(new_n475), .C2(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n461), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n481), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n492), .A2(KEYINPUT69), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n492), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n503), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT70), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n511), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n503), .A2(new_n504), .A3(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n504), .A2(KEYINPUT72), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT73), .B(G51), .Z(new_n531));
  NAND3_X1  g106(.A1(new_n501), .A2(KEYINPUT71), .A3(new_n502), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  AND2_X1   g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n530), .A2(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n525), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n526), .B1(new_n525), .B2(new_n539), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n512), .ZN(new_n546));
  INV_X1    g121(.A(new_n505), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n530), .A2(G52), .B1(new_n547), .B2(G90), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n530), .A2(G43), .B1(new_n547), .B2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n532), .A2(new_n536), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n547), .A2(new_n563), .A3(G91), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n505), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n510), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n510), .B2(new_n567), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n564), .A2(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n512), .B1(new_n571), .B2(KEYINPUT77), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n572), .B1(KEYINPUT77), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n546), .A2(new_n548), .ZN(G301));
  INV_X1    g150(.A(G166), .ZN(G303));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n552), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n578), .A2(KEYINPUT78), .A3(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n532), .B2(new_n536), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n512), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n510), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n547), .A2(G87), .B1(G49), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G61), .B1(new_n534), .B2(new_n535), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(KEYINPUT79), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n503), .A2(new_n591), .A3(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n512), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n503), .A2(new_n504), .A3(G86), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n512), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n530), .A2(G47), .B1(new_n547), .B2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  AND3_X1   g177(.A1(new_n503), .A2(new_n504), .A3(G92), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n530), .A2(G54), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n503), .A2(G66), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G171), .B2(new_n610), .ZN(G284));
  OAI21_X1  g187(.A(new_n611), .B1(G171), .B2(new_n610), .ZN(G321));
  NOR2_X1   g188(.A1(G286), .A2(new_n610), .ZN(new_n614));
  XOR2_X1   g189(.A(G299), .B(KEYINPUT80), .Z(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n610), .B2(new_n615), .ZN(G297));
  XNOR2_X1  g191(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g192(.A(new_n609), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n556), .A2(new_n610), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n609), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n462), .A2(new_n468), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n477), .A2(G135), .B1(G123), .B2(new_n481), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n632), .A2(new_n461), .A3(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n461), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n629), .A2(new_n630), .A3(new_n638), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n640));
  INV_X1    g215(.A(G1341), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT83), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT84), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n646), .A2(new_n650), .A3(KEYINPUT14), .A4(new_n647), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n641), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G1348), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n641), .A3(new_n651), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n649), .A2(new_n641), .A3(new_n651), .ZN(new_n657));
  OAI21_X1  g232(.A(G1348), .B1(new_n657), .B2(new_n652), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n662), .B1(new_n656), .B2(new_n658), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n640), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n665), .ZN(new_n667));
  NAND4_X1  g242(.A1(new_n667), .A2(KEYINPUT85), .A3(G14), .A4(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n628), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n637), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n695), .B(new_n694), .S(new_n687), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n693), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n693), .B2(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT86), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n703), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n684), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(new_n683), .A3(new_n704), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G20), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT23), .Z(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G299), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1956), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  INV_X1    g293(.A(G127), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n476), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n461), .B1(new_n720), .B2(KEYINPUT89), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT89), .B2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n723));
  NAND2_X1  g298(.A1(G103), .A2(G2104), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G2105), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n477), .A2(G139), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G33), .B(new_n728), .S(G29), .Z(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G2072), .Z(new_n730));
  NOR2_X1   g305(.A1(G29), .A2(G35), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G162), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2090), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G1996), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n468), .A2(G105), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n741), .B(new_n742), .C1(G141), .C2(new_n477), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n481), .A2(G129), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n738), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT27), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n717), .B(new_n736), .C1(new_n737), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n738), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n477), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n481), .A2(G128), .ZN(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n738), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n738), .B1(new_n763), .B2(G28), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n763), .B2(G28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(KEYINPUT92), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n769), .B2(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT24), .B2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n463), .A2(new_n465), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n461), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n771), .B1(new_n774), .B2(new_n738), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n768), .B1(new_n738), .B2(new_n636), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n761), .B(new_n778), .C1(new_n749), .C2(new_n737), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n712), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n618), .B2(new_n712), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1348), .ZN(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G19), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n557), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT88), .B(G1341), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n779), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G286), .A2(G16), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n712), .A2(G21), .ZN(new_n789));
  INV_X1    g364(.A(G1966), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n788), .A2(new_n789), .B1(KEYINPUT91), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  NOR2_X1   g368(.A1(G5), .A2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G301), .B2(new_n712), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n738), .A2(G27), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT94), .Z(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n738), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n750), .A2(new_n787), .A3(new_n793), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n712), .A2(G23), .ZN(new_n805));
  INV_X1    g380(.A(G288), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n712), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n712), .A2(G22), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G166), .B2(new_n712), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1971), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n712), .A2(G6), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n597), .B2(new_n712), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT32), .B(G1981), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n812), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n809), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n712), .A2(G24), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n600), .A2(new_n601), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n712), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1986), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n481), .A2(G119), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n461), .A2(G107), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(G131), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n826), .B1(new_n827), .B2(new_n828), .C1(new_n829), .C2(new_n470), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT87), .ZN(new_n831));
  MUX2_X1   g406(.A(G25), .B(new_n831), .S(G29), .Z(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n825), .B(new_n834), .C1(new_n819), .C2(KEYINPUT34), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT36), .B1(new_n821), .B2(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n821), .A2(new_n835), .A3(KEYINPUT36), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n804), .B1(new_n836), .B2(new_n837), .ZN(G311));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  XNOR2_X1  g414(.A(G311), .B(new_n839), .ZN(G150));
  AOI22_X1  g415(.A1(new_n530), .A2(G55), .B1(new_n547), .B2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n537), .A2(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g419(.A(KEYINPUT97), .B(new_n841), .C1(new_n844), .C2(new_n512), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n846));
  INV_X1    g421(.A(new_n841), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n512), .B1(new_n842), .B2(new_n843), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n557), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n556), .A2(new_n847), .A3(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n619), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n845), .A2(new_n849), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(G162), .B(G160), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT98), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(new_n636), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n636), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n481), .A2(G126), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n493), .A2(new_n495), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n872));
  INV_X1    g447(.A(new_n491), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n490), .B1(new_n462), .B2(new_n487), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n489), .A2(KEYINPUT99), .A3(new_n491), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n758), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(new_n831), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n728), .B(new_n746), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n481), .A2(G130), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n461), .A2(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n881), .B1(new_n882), .B2(new_n883), .C1(new_n884), .C2(new_n470), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n626), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n880), .A2(new_n886), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n886), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n880), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n878), .B(new_n831), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n868), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n892), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n895), .B(new_n896), .C1(new_n867), .C2(new_n866), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g475(.A1(new_n850), .A2(new_n851), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n622), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n609), .B(G299), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(KEYINPUT41), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT102), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G290), .A2(G288), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(G290), .A2(G288), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n597), .B(G303), .ZN(new_n914));
  OR4_X1    g489(.A1(KEYINPUT101), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT101), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n913), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n911), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n904), .A2(KEYINPUT102), .A3(new_n909), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n910), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n910), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(G868), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G868), .B2(new_n859), .ZN(G295));
  OAI21_X1  g502(.A(new_n926), .B1(G868), .B2(new_n859), .ZN(G331));
  AND3_X1   g503(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n523), .B1(new_n518), .B2(new_n520), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n530), .A2(new_n531), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n537), .A2(new_n538), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT75), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(G171), .A2(new_n540), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(G301), .B1(new_n541), .B2(new_n542), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n852), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(new_n903), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n852), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT103), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n852), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n915), .A2(new_n920), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n936), .B(new_n937), .C1(new_n850), .C2(new_n851), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n908), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n947), .A3(new_n944), .ZN(new_n951));
  MUX2_X1   g526(.A(new_n905), .B(KEYINPUT41), .S(new_n903), .Z(new_n952));
  AOI22_X1  g527(.A1(new_n951), .A2(new_n952), .B1(new_n941), .B2(new_n940), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n950), .B(new_n898), .C1(new_n953), .C2(new_n946), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n938), .A2(new_n852), .A3(new_n943), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n943), .B1(new_n938), .B2(new_n852), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n959), .A2(new_n940), .B1(new_n948), .B2(new_n908), .ZN(new_n960));
  AOI21_X1  g535(.A(G37), .B1(new_n960), .B2(new_n946), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n946), .B1(new_n945), .B2(new_n949), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT44), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n951), .A2(new_n952), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n940), .A2(new_n941), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n921), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n961), .A3(new_n955), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n950), .A2(new_n898), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT43), .B1(new_n970), .B2(new_n962), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n965), .B1(new_n973), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n877), .B2(G1384), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT104), .B(G40), .Z(new_n977));
  NOR3_X1   g552(.A1(new_n466), .A2(new_n472), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n757), .B(new_n760), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n983), .A2(KEYINPUT105), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(KEYINPUT105), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n746), .B(G1996), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n984), .A2(new_n985), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n833), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n831), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n758), .A2(new_n760), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n980), .A2(new_n737), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n982), .A2(new_n747), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n993), .A2(new_n994), .B1(new_n980), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  AND2_X1   g575(.A1(new_n831), .A2(new_n988), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n980), .B1(new_n1001), .B2(new_n989), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n987), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  AOI211_X1 g580(.A(new_n992), .B(new_n1000), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT106), .B(G8), .Z(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n935), .A2(new_n540), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT122), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n935), .A2(new_n540), .A3(KEYINPUT122), .A4(new_n1008), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT69), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n873), .A2(new_n874), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(new_n871), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n492), .A2(KEYINPUT69), .A3(new_n496), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(KEYINPUT45), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n976), .A2(new_n978), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n790), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n489), .A2(KEYINPUT99), .A3(new_n491), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT99), .B1(new_n489), .B2(new_n491), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n496), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n1017), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT114), .B(G2084), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1023), .A2(new_n978), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1013), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1021), .A2(new_n1011), .A3(new_n1030), .A4(new_n1012), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(KEYINPUT51), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1007), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1011), .A2(new_n1036), .A3(new_n1012), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1033), .A2(KEYINPUT51), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1032), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1022), .A2(new_n975), .ZN(new_n1045));
  INV_X1    g620(.A(G2078), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1026), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n978), .A4(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1023), .A2(new_n978), .A3(new_n1028), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1048), .A2(new_n1049), .B1(new_n1050), .B2(new_n797), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(KEYINPUT53), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1020), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G301), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G166), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT55), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n499), .A2(new_n1058), .A3(new_n1027), .A4(new_n1017), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1016), .A2(new_n1027), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT113), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1027), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n979), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n875), .A2(new_n876), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1384), .B1(new_n1067), .B2(new_n496), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT112), .B(new_n978), .C1(new_n1068), .C2(new_n1027), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n979), .B1(new_n1068), .B2(KEYINPUT45), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1971), .B1(new_n1071), .B2(new_n1045), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1057), .B1(new_n1074), .B2(new_n1008), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  INV_X1    g651(.A(G1981), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n589), .A2(KEYINPUT79), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n592), .A2(new_n1078), .A3(new_n587), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n596), .B1(new_n1079), .B2(G651), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT108), .B(G86), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n547), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1077), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NOR4_X1   g658(.A1(new_n593), .A2(G1981), .A3(new_n594), .A4(new_n596), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT109), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT109), .B(new_n1076), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1026), .A2(new_n1017), .A3(new_n978), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1008), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(KEYINPUT49), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT52), .B(G1976), .C1(new_n583), .C2(new_n585), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT78), .B1(new_n578), .B2(G651), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n581), .A2(new_n580), .A3(new_n512), .ZN(new_n1096));
  OAI211_X1 g671(.A(G1976), .B(new_n585), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(new_n1008), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(KEYINPUT107), .A2(KEYINPUT52), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1090), .A2(new_n1008), .A3(new_n1097), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1089), .A2(new_n1093), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1066), .A2(new_n1023), .A3(new_n978), .A4(new_n1028), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1057), .C1(new_n1104), .C2(new_n1072), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1075), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1040), .A2(new_n1044), .A3(new_n1054), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1007), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1105), .B(new_n1103), .C1(new_n1110), .C2(new_n1057), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1035), .A2(G168), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1109), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1104), .A2(new_n1072), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1055), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1057), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1084), .B(KEYINPUT110), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT111), .Z(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1091), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1105), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(new_n1124), .B1(new_n1125), .B2(new_n1103), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1108), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  OAI21_X1  g703(.A(G299), .B1(KEYINPUT116), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(KEYINPUT116), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT117), .Z(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1129), .B(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1071), .A2(new_n1045), .A3(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1062), .A2(new_n1069), .A3(new_n1065), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n716), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1137), .B2(new_n716), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1090), .A2(G2067), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1050), .B2(new_n654), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n609), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT118), .Z(new_n1145));
  NAND2_X1  g720(.A1(new_n1137), .A2(new_n716), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT115), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1137), .A2(new_n1138), .A3(new_n716), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1133), .B1(new_n1149), .B2(new_n1135), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1141), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1141), .A2(KEYINPUT61), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT120), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1133), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT61), .A4(new_n1141), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1143), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT121), .B(new_n618), .C1(new_n1143), .C2(KEYINPUT60), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1050), .A2(new_n654), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1142), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(KEYINPUT60), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n609), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1071), .A2(new_n737), .A3(new_n1045), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT58), .B(G1341), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1090), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1170), .A2(KEYINPUT119), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT119), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n557), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT59), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1154), .A2(new_n1155), .B1(new_n1149), .B2(new_n1136), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1169), .B(new_n1176), .C1(new_n1177), .C2(KEYINPUT61), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1151), .B1(new_n1159), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1050), .A2(new_n797), .ZN(new_n1182));
  INV_X1    g757(.A(G40), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n774), .A2(new_n1183), .A3(new_n1052), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n976), .A2(new_n1047), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(G171), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1180), .B1(new_n1187), .B2(new_n1054), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1107), .A2(new_n1188), .A3(new_n1043), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1051), .A2(G301), .A3(new_n1053), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT54), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1186), .A2(KEYINPUT124), .ZN(new_n1192));
  AOI21_X1  g767(.A(G301), .B1(new_n1186), .B2(KEYINPUT124), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT125), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1038), .A2(new_n1111), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1191), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1196), .A2(new_n1199), .A3(new_n1200), .A4(new_n1188), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1127), .B1(new_n1179), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n823), .B(G1986), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1003), .B1(new_n981), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1006), .B1(new_n1203), .B2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g781(.A1(G227), .A2(new_n459), .ZN(new_n1208));
  AND3_X1   g782(.A1(new_n707), .A2(new_n709), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n669), .A2(new_n899), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g784(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g785(.A(KEYINPUT127), .B1(new_n972), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  AOI211_X1 g787(.A(new_n1213), .B(new_n1210), .C1(new_n969), .C2(new_n971), .ZN(new_n1214));
  NOR2_X1   g788(.A1(new_n1212), .A2(new_n1214), .ZN(G308));
  NOR2_X1   g789(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n955), .B1(new_n961), .B2(new_n963), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1211), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(new_n1213), .ZN(new_n1219));
  NAND3_X1  g793(.A1(new_n972), .A2(KEYINPUT127), .A3(new_n1211), .ZN(new_n1220));
  NAND2_X1  g794(.A1(new_n1219), .A2(new_n1220), .ZN(G225));
endmodule


