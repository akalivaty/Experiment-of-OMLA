

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769;

  NOR2_X2 U376 ( .A1(n545), .A2(n524), .ZN(n727) );
  XNOR2_X1 U377 ( .A(n419), .B(G953), .ZN(n474) );
  BUF_X2 U378 ( .A(n474), .Z(n671) );
  NOR2_X2 U379 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X2 U380 ( .A(n366), .B(n430), .ZN(n530) );
  NAND2_X2 U381 ( .A1(n427), .A2(n609), .ZN(n366) );
  XNOR2_X1 U382 ( .A(G902), .B(KEYINPUT87), .ZN(n426) );
  BUF_X1 U383 ( .A(n690), .Z(n697) );
  XNOR2_X1 U384 ( .A(n669), .B(G146), .ZN(n367) );
  XNOR2_X1 U385 ( .A(G116), .B(G113), .ZN(n401) );
  NAND2_X1 U386 ( .A1(n379), .A2(n511), .ZN(n578) );
  OR2_X1 U387 ( .A1(n575), .A2(n357), .ZN(n378) );
  NOR2_X1 U388 ( .A1(n731), .A2(n592), .ZN(n583) );
  XNOR2_X1 U389 ( .A(n389), .B(n365), .ZN(n575) );
  XNOR2_X1 U390 ( .A(n582), .B(n581), .ZN(n731) );
  NAND2_X1 U391 ( .A1(n386), .A2(n385), .ZN(n381) );
  XNOR2_X1 U392 ( .A(n392), .B(n391), .ZN(n520) );
  XNOR2_X1 U393 ( .A(n499), .B(n498), .ZN(n513) );
  AND2_X1 U394 ( .A1(n691), .A2(n494), .ZN(n499) );
  XNOR2_X1 U395 ( .A(n395), .B(KEYINPUT20), .ZN(n495) );
  XNOR2_X1 U396 ( .A(n402), .B(n401), .ZN(n501) );
  XNOR2_X1 U397 ( .A(n380), .B(G119), .ZN(n402) );
  XNOR2_X1 U398 ( .A(G107), .B(G104), .ZN(n414) );
  INV_X2 U399 ( .A(KEYINPUT64), .ZN(n419) );
  INV_X2 U400 ( .A(KEYINPUT3), .ZN(n380) );
  XNOR2_X1 U401 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n412) );
  XNOR2_X2 U402 ( .A(KEYINPUT109), .B(n537), .ZN(n722) );
  XNOR2_X2 U403 ( .A(n570), .B(n569), .ZN(n572) );
  XNOR2_X2 U404 ( .A(n444), .B(n443), .ZN(n481) );
  XNOR2_X2 U405 ( .A(n530), .B(KEYINPUT38), .ZN(n725) );
  XNOR2_X2 U406 ( .A(n521), .B(KEYINPUT79), .ZN(n531) );
  BUF_X1 U407 ( .A(n739), .Z(n353) );
  XNOR2_X1 U408 ( .A(n534), .B(KEYINPUT1), .ZN(n739) );
  AND2_X1 U409 ( .A1(n578), .A2(n658), .ZN(n586) );
  XNOR2_X1 U410 ( .A(n398), .B(n438), .ZN(n515) );
  INV_X1 U411 ( .A(KEYINPUT91), .ZN(n438) );
  INV_X1 U412 ( .A(KEYINPUT106), .ZN(n397) );
  INV_X1 U413 ( .A(G237), .ZN(n428) );
  XNOR2_X1 U414 ( .A(n472), .B(G137), .ZN(n390) );
  XNOR2_X1 U415 ( .A(n608), .B(n607), .ZN(n623) );
  INV_X1 U416 ( .A(KEYINPUT45), .ZN(n607) );
  XOR2_X1 U417 ( .A(G131), .B(G140), .Z(n476) );
  XNOR2_X1 U418 ( .A(G146), .B(G125), .ZN(n465) );
  XNOR2_X1 U419 ( .A(n478), .B(G469), .ZN(n479) );
  XNOR2_X1 U420 ( .A(n500), .B(n400), .ZN(n399) );
  XNOR2_X1 U421 ( .A(G131), .B(G101), .ZN(n500) );
  XNOR2_X1 U422 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n400) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n502) );
  XNOR2_X1 U424 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U425 ( .A(G140), .ZN(n489) );
  XNOR2_X1 U426 ( .A(G128), .B(G119), .ZN(n490) );
  XNOR2_X1 U427 ( .A(n486), .B(KEYINPUT93), .ZN(n487) );
  INV_X1 U428 ( .A(KEYINPUT92), .ZN(n486) );
  XNOR2_X1 U429 ( .A(n538), .B(n539), .ZN(n752) );
  OR2_X1 U430 ( .A1(n643), .A2(G902), .ZN(n506) );
  NAND2_X1 U431 ( .A1(n382), .A2(n381), .ZN(n389) );
  AND2_X1 U432 ( .A1(n388), .A2(n383), .ZN(n382) );
  NAND2_X1 U433 ( .A1(n733), .A2(KEYINPUT70), .ZN(n403) );
  NAND2_X1 U434 ( .A1(n442), .A2(KEYINPUT0), .ZN(n387) );
  XNOR2_X1 U435 ( .A(G143), .B(G113), .ZN(n454) );
  NOR2_X1 U436 ( .A1(n612), .A2(n611), .ZN(n615) );
  XNOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n418) );
  XNOR2_X1 U438 ( .A(n435), .B(KEYINPUT77), .ZN(n436) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n435) );
  NOR2_X1 U440 ( .A1(n518), .A2(n355), .ZN(n525) );
  XNOR2_X1 U441 ( .A(n396), .B(n397), .ZN(n516) );
  OR2_X1 U442 ( .A1(n737), .A2(n432), .ZN(n392) );
  INV_X1 U443 ( .A(KEYINPUT30), .ZN(n391) );
  NAND2_X1 U444 ( .A1(n406), .A2(n404), .ZN(n533) );
  NAND2_X1 U445 ( .A1(n410), .A2(n405), .ZN(n404) );
  AND2_X1 U446 ( .A1(n407), .A2(n409), .ZN(n406) );
  NOR2_X1 U447 ( .A1(n734), .A2(n403), .ZN(n405) );
  INV_X1 U448 ( .A(G902), .ZN(n494) );
  NAND2_X1 U449 ( .A1(n542), .A2(KEYINPUT0), .ZN(n388) );
  XNOR2_X1 U450 ( .A(G116), .B(G107), .ZN(n447) );
  XNOR2_X1 U451 ( .A(n376), .B(n477), .ZN(n375) );
  XNOR2_X1 U452 ( .A(n475), .B(n377), .ZN(n376) );
  XNOR2_X1 U453 ( .A(n367), .B(n505), .ZN(n643) );
  XNOR2_X1 U454 ( .A(n501), .B(n399), .ZN(n504) );
  XNOR2_X1 U455 ( .A(n393), .B(n488), .ZN(n492) );
  XNOR2_X1 U456 ( .A(n491), .B(n487), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n368), .B(n540), .ZN(n767) );
  NOR2_X1 U458 ( .A1(n543), .A2(n752), .ZN(n368) );
  INV_X1 U459 ( .A(KEYINPUT40), .ZN(n369) );
  NOR2_X1 U460 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U461 ( .A(n373), .B(n372), .ZN(n585) );
  INV_X1 U462 ( .A(KEYINPUT35), .ZN(n372) );
  XNOR2_X1 U463 ( .A(n583), .B(KEYINPUT34), .ZN(n374) );
  NOR2_X1 U464 ( .A1(n543), .A2(n542), .ZN(n711) );
  AND2_X1 U465 ( .A1(n572), .A2(n571), .ZN(n354) );
  XOR2_X1 U466 ( .A(KEYINPUT107), .B(n517), .Z(n355) );
  XNOR2_X1 U467 ( .A(n465), .B(n464), .ZN(n488) );
  AND2_X1 U468 ( .A1(n533), .A2(n371), .ZN(n356) );
  OR2_X1 U469 ( .A1(n577), .A2(n579), .ZN(n357) );
  AND2_X1 U470 ( .A1(n566), .A2(n720), .ZN(n358) );
  OR2_X1 U471 ( .A1(n734), .A2(n411), .ZN(n359) );
  AND2_X1 U472 ( .A1(n567), .A2(n358), .ZN(n360) );
  INV_X1 U473 ( .A(n733), .ZN(n411) );
  AND2_X1 U474 ( .A1(n571), .A2(n721), .ZN(n361) );
  AND2_X1 U475 ( .A1(n625), .A2(KEYINPUT81), .ZN(n362) );
  AND2_X1 U476 ( .A1(n354), .A2(n362), .ZN(n363) );
  AND2_X1 U477 ( .A1(n388), .A2(n387), .ZN(n364) );
  XOR2_X1 U478 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n365) );
  XNOR2_X1 U479 ( .A(n532), .B(KEYINPUT39), .ZN(n573) );
  XNOR2_X2 U480 ( .A(n434), .B(n433), .ZN(n542) );
  NAND2_X1 U481 ( .A1(n536), .A2(n535), .ZN(n543) );
  AND2_X2 U482 ( .A1(n572), .A2(n361), .ZN(n666) );
  AND2_X2 U483 ( .A1(n623), .A2(n666), .ZN(n619) );
  NAND2_X1 U484 ( .A1(n585), .A2(n586), .ZN(n589) );
  NOR2_X1 U485 ( .A1(n652), .A2(G902), .ZN(n480) );
  XNOR2_X1 U486 ( .A(n375), .B(n367), .ZN(n652) );
  NOR2_X2 U487 ( .A1(n768), .A2(n767), .ZN(n541) );
  XNOR2_X2 U488 ( .A(n370), .B(n369), .ZN(n768) );
  NAND2_X1 U489 ( .A1(n573), .A2(n713), .ZN(n370) );
  XNOR2_X2 U490 ( .A(n506), .B(n641), .ZN(n737) );
  AND2_X1 U491 ( .A1(n576), .A2(n737), .ZN(n511) );
  NOR2_X1 U492 ( .A1(n595), .A2(n371), .ZN(n597) );
  INV_X1 U493 ( .A(n737), .ZN(n371) );
  INV_X1 U494 ( .A(n585), .ZN(n765) );
  NAND2_X1 U495 ( .A1(n374), .A2(n584), .ZN(n373) );
  INV_X1 U496 ( .A(n476), .ZN(n377) );
  XNOR2_X2 U497 ( .A(n473), .B(n390), .ZN(n669) );
  XNOR2_X2 U498 ( .A(n378), .B(KEYINPUT32), .ZN(n658) );
  XNOR2_X1 U499 ( .A(n510), .B(KEYINPUT104), .ZN(n379) );
  NAND2_X1 U500 ( .A1(n364), .A2(n381), .ZN(n592) );
  NOR2_X1 U501 ( .A1(n471), .A2(n384), .ZN(n383) );
  INV_X1 U502 ( .A(n387), .ZN(n384) );
  NOR2_X1 U503 ( .A1(n442), .A2(KEYINPUT0), .ZN(n385) );
  INV_X1 U504 ( .A(n542), .ZN(n386) );
  NOR2_X2 U505 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X2 U506 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n472) );
  XNOR2_X2 U507 ( .A(n449), .B(G134), .ZN(n473) );
  XNOR2_X2 U508 ( .A(G143), .B(G128), .ZN(n449) );
  XNOR2_X2 U509 ( .A(n394), .B(n469), .ZN(n733) );
  NAND2_X1 U510 ( .A1(n495), .A2(G221), .ZN(n394) );
  NAND2_X1 U511 ( .A1(n609), .A2(G234), .ZN(n395) );
  NOR2_X2 U512 ( .A1(n515), .A2(n671), .ZN(n396) );
  NAND2_X1 U513 ( .A1(n440), .A2(G902), .ZN(n398) );
  NAND2_X1 U514 ( .A1(n525), .A2(n408), .ZN(n409) );
  NAND2_X1 U515 ( .A1(n359), .A2(n408), .ZN(n407) );
  INV_X1 U516 ( .A(KEYINPUT70), .ZN(n408) );
  INV_X1 U517 ( .A(n525), .ZN(n410) );
  XNOR2_X2 U518 ( .A(n426), .B(n425), .ZN(n609) );
  INV_X1 U519 ( .A(KEYINPUT48), .ZN(n569) );
  XNOR2_X1 U520 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n581) );
  BUF_X1 U521 ( .A(n666), .Z(n670) );
  BUF_X1 U522 ( .A(n530), .Z(n562) );
  XNOR2_X1 U523 ( .A(n412), .B(G122), .ZN(n413) );
  XNOR2_X1 U524 ( .A(n501), .B(n413), .ZN(n417) );
  XNOR2_X1 U525 ( .A(n414), .B(G110), .ZN(n416) );
  XNOR2_X1 U526 ( .A(G101), .B(KEYINPUT78), .ZN(n415) );
  XNOR2_X1 U527 ( .A(n416), .B(n415), .ZN(n477) );
  XNOR2_X1 U528 ( .A(n417), .B(n477), .ZN(n686) );
  XNOR2_X1 U529 ( .A(n449), .B(n418), .ZN(n421) );
  NAND2_X1 U530 ( .A1(n671), .A2(G224), .ZN(n420) );
  XNOR2_X1 U531 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X1 U532 ( .A(n472), .B(n465), .ZN(n422) );
  XNOR2_X1 U533 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U534 ( .A(n686), .B(n424), .ZN(n630) );
  INV_X1 U535 ( .A(n630), .ZN(n427) );
  INV_X1 U536 ( .A(KEYINPUT15), .ZN(n425) );
  NAND2_X1 U537 ( .A1(n494), .A2(n428), .ZN(n431) );
  NAND2_X1 U538 ( .A1(n431), .A2(G210), .ZN(n429) );
  XNOR2_X1 U539 ( .A(n429), .B(KEYINPUT80), .ZN(n430) );
  NAND2_X1 U540 ( .A1(n431), .A2(G214), .ZN(n724) );
  INV_X1 U541 ( .A(n724), .ZN(n432) );
  OR2_X2 U542 ( .A1(n530), .A2(n432), .ZN(n434) );
  XNOR2_X1 U543 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n433) );
  XOR2_X1 U544 ( .A(KEYINPUT88), .B(KEYINPUT14), .Z(n437) );
  XNOR2_X1 U545 ( .A(n437), .B(n436), .ZN(n440) );
  XNOR2_X1 U546 ( .A(G898), .B(KEYINPUT89), .ZN(n683) );
  NAND2_X1 U547 ( .A1(n683), .A2(G953), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n439), .B(KEYINPUT90), .ZN(n687) );
  NOR2_X1 U549 ( .A1(n515), .A2(n687), .ZN(n441) );
  NAND2_X1 U550 ( .A1(G952), .A2(n440), .ZN(n751) );
  NOR2_X1 U551 ( .A1(n751), .A2(G953), .ZN(n518) );
  NOR2_X1 U552 ( .A1(n441), .A2(n518), .ZN(n442) );
  XOR2_X1 U553 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n446) );
  NAND2_X1 U554 ( .A1(n474), .A2(G234), .ZN(n444) );
  INV_X1 U555 ( .A(KEYINPUT8), .ZN(n443) );
  NAND2_X1 U556 ( .A1(G217), .A2(n481), .ZN(n445) );
  XNOR2_X1 U557 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U558 ( .A(KEYINPUT7), .B(G122), .Z(n448) );
  XNOR2_X1 U559 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U560 ( .A(n473), .B(n450), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n699) );
  NAND2_X1 U562 ( .A1(n699), .A2(n494), .ZN(n453) );
  XNOR2_X1 U563 ( .A(n453), .B(G478), .ZN(n545) );
  XOR2_X1 U564 ( .A(G122), .B(G104), .Z(n455) );
  XNOR2_X1 U565 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U566 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n457) );
  XNOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT11), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n463) );
  XOR2_X1 U570 ( .A(KEYINPUT99), .B(KEYINPUT102), .Z(n461) );
  NAND2_X1 U571 ( .A1(G214), .A2(n502), .ZN(n460) );
  XOR2_X1 U572 ( .A(n461), .B(n460), .Z(n462) );
  XNOR2_X1 U573 ( .A(n463), .B(n462), .ZN(n466) );
  INV_X1 U574 ( .A(KEYINPUT10), .ZN(n464) );
  XNOR2_X1 U575 ( .A(n476), .B(n488), .ZN(n667) );
  XNOR2_X1 U576 ( .A(n466), .B(n667), .ZN(n660) );
  NAND2_X1 U577 ( .A1(n660), .A2(n494), .ZN(n468) );
  XOR2_X1 U578 ( .A(KEYINPUT13), .B(G475), .Z(n467) );
  XNOR2_X1 U579 ( .A(n468), .B(n467), .ZN(n524) );
  INV_X1 U580 ( .A(KEYINPUT21), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n733), .B(KEYINPUT95), .ZN(n512) );
  INV_X1 U582 ( .A(n512), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n727), .A2(n470), .ZN(n471) );
  NAND2_X1 U584 ( .A1(n671), .A2(G227), .ZN(n475) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n478) );
  XNOR2_X2 U586 ( .A(n480), .B(n479), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n481), .A2(G221), .ZN(n485) );
  XOR2_X1 U588 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n483) );
  XNOR2_X1 U589 ( .A(G137), .B(G110), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n485), .B(n484), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n493), .B(n492), .ZN(n691) );
  NAND2_X1 U593 ( .A1(n495), .A2(G217), .ZN(n497) );
  XNOR2_X1 U594 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n496) );
  XOR2_X1 U595 ( .A(n497), .B(n496), .Z(n498) );
  INV_X1 U596 ( .A(n513), .ZN(n734) );
  INV_X1 U597 ( .A(n734), .ZN(n576) );
  NOR2_X1 U598 ( .A1(n353), .A2(n576), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n502), .A2(G210), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U601 ( .A(G472), .ZN(n641) );
  XNOR2_X1 U602 ( .A(n737), .B(KEYINPUT6), .ZN(n579) );
  INV_X1 U603 ( .A(n579), .ZN(n507) );
  NAND2_X1 U604 ( .A1(n508), .A2(n507), .ZN(n509) );
  OR2_X1 U605 ( .A1(n575), .A2(n509), .ZN(n602) );
  XNOR2_X1 U606 ( .A(n602), .B(G101), .ZN(G3) );
  NOR2_X1 U607 ( .A1(n575), .A2(n353), .ZN(n510) );
  XNOR2_X1 U608 ( .A(n578), .B(G110), .ZN(G12) );
  XNOR2_X2 U609 ( .A(n514), .B(KEYINPUT68), .ZN(n738) );
  NAND2_X1 U610 ( .A1(n738), .A2(n534), .ZN(n595) );
  NOR2_X1 U611 ( .A1(G900), .A2(n516), .ZN(n517) );
  NOR2_X1 U612 ( .A1(n595), .A2(n525), .ZN(n519) );
  NAND2_X1 U613 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U614 ( .A1(n545), .A2(n524), .ZN(n522) );
  XNOR2_X1 U615 ( .A(KEYINPUT105), .B(n522), .ZN(n584) );
  NAND2_X1 U616 ( .A1(n531), .A2(n584), .ZN(n523) );
  OR2_X1 U617 ( .A1(n562), .A2(n523), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(G143), .ZN(G45) );
  INV_X1 U619 ( .A(n524), .ZN(n544) );
  OR2_X1 U620 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U621 ( .A1(n579), .A2(n533), .ZN(n526) );
  NOR2_X1 U622 ( .A1(n546), .A2(n526), .ZN(n527) );
  NAND2_X1 U623 ( .A1(n527), .A2(n724), .ZN(n563) );
  OR2_X1 U624 ( .A1(n563), .A2(n353), .ZN(n528) );
  XNOR2_X1 U625 ( .A(KEYINPUT43), .B(n528), .ZN(n529) );
  NAND2_X1 U626 ( .A1(n529), .A2(n562), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(G140), .ZN(G42) );
  NAND2_X1 U628 ( .A1(n531), .A2(n725), .ZN(n532) );
  INV_X1 U629 ( .A(n546), .ZN(n713) );
  XNOR2_X1 U630 ( .A(n356), .B(KEYINPUT28), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n534), .B(KEYINPUT108), .ZN(n535) );
  XOR2_X1 U632 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n539) );
  NAND2_X1 U633 ( .A1(n725), .A2(n724), .ZN(n537) );
  NAND2_X1 U634 ( .A1(n722), .A2(n727), .ZN(n538) );
  XOR2_X1 U635 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n540) );
  XNOR2_X1 U636 ( .A(n541), .B(KEYINPUT46), .ZN(n568) );
  AND2_X1 U637 ( .A1(n545), .A2(n544), .ZN(n716) );
  INV_X1 U638 ( .A(n716), .ZN(n547) );
  NAND2_X1 U639 ( .A1(n547), .A2(n546), .ZN(n723) );
  INV_X1 U640 ( .A(n723), .ZN(n551) );
  NOR2_X1 U641 ( .A1(n551), .A2(KEYINPUT69), .ZN(n548) );
  NAND2_X1 U642 ( .A1(n711), .A2(n548), .ZN(n549) );
  INV_X1 U643 ( .A(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n549), .A2(n557), .ZN(n556) );
  AND2_X1 U645 ( .A1(n551), .A2(KEYINPUT82), .ZN(n553) );
  NOR2_X1 U646 ( .A1(n557), .A2(KEYINPUT69), .ZN(n550) );
  NOR2_X1 U647 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U648 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U649 ( .A1(n711), .A2(n554), .ZN(n555) );
  NAND2_X1 U650 ( .A1(n556), .A2(n555), .ZN(n567) );
  NOR2_X1 U651 ( .A1(n557), .A2(n723), .ZN(n558) );
  NOR2_X1 U652 ( .A1(KEYINPUT82), .A2(n558), .ZN(n561) );
  INV_X1 U653 ( .A(n559), .ZN(n560) );
  NOR2_X1 U654 ( .A1(n561), .A2(n560), .ZN(n566) );
  XNOR2_X1 U655 ( .A(n564), .B(KEYINPUT36), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n565), .A2(n353), .ZN(n720) );
  NAND2_X1 U657 ( .A1(n568), .A2(n360), .ZN(n570) );
  BUF_X1 U658 ( .A(n573), .Z(n574) );
  NAND2_X1 U659 ( .A1(n574), .A2(n716), .ZN(n721) );
  NAND2_X1 U660 ( .A1(n353), .A2(n576), .ZN(n577) );
  NAND2_X1 U661 ( .A1(n739), .A2(n738), .ZN(n590) );
  INV_X1 U662 ( .A(n590), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n587), .A2(KEYINPUT74), .ZN(n588) );
  XNOR2_X1 U666 ( .A(n589), .B(n588), .ZN(n606) );
  NOR2_X1 U667 ( .A1(n737), .A2(n590), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT98), .B(n591), .ZN(n743) );
  INV_X1 U669 ( .A(n592), .ZN(n596) );
  AND2_X1 U670 ( .A1(n743), .A2(n596), .ZN(n594) );
  INV_X1 U671 ( .A(KEYINPUT31), .ZN(n593) );
  XNOR2_X1 U672 ( .A(n594), .B(n593), .ZN(n717) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT97), .ZN(n706) );
  OR2_X1 U675 ( .A1(n717), .A2(n706), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n599), .A2(n723), .ZN(n604) );
  INV_X1 U677 ( .A(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n600), .A2(KEYINPUT44), .ZN(n601) );
  AND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U681 ( .A(n609), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n619), .A2(n613), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n610), .A2(KEYINPUT83), .ZN(n617) );
  NAND2_X1 U684 ( .A1(n623), .A2(n666), .ZN(n612) );
  OR2_X1 U685 ( .A1(KEYINPUT83), .A2(n609), .ZN(n611) );
  AND2_X1 U686 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT66), .ZN(n628) );
  INV_X1 U690 ( .A(n619), .ZN(n620) );
  INV_X1 U691 ( .A(n620), .ZN(n757) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n621), .A2(KEYINPUT81), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n757), .A2(n622), .ZN(n627) );
  BUF_X1 U695 ( .A(n623), .Z(n624) );
  NAND2_X1 U696 ( .A1(n721), .A2(KEYINPUT2), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n624), .A2(n363), .ZN(n626) );
  AND2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n756) );
  NAND2_X2 U699 ( .A1(n628), .A2(n756), .ZN(n648) );
  INV_X1 U700 ( .A(G210), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n648), .A2(n629), .ZN(n635) );
  BUF_X1 U702 ( .A(n630), .Z(n631) );
  XNOR2_X1 U703 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n632) );
  XOR2_X1 U704 ( .A(n632), .B(KEYINPUT55), .Z(n633) );
  XNOR2_X1 U705 ( .A(n631), .B(n633), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n638) );
  INV_X1 U707 ( .A(n671), .ZN(n637) );
  INV_X1 U708 ( .A(G952), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n695) );
  NAND2_X1 U710 ( .A1(n638), .A2(n695), .ZN(n640) );
  INV_X1 U711 ( .A(KEYINPUT56), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(G51) );
  NOR2_X1 U713 ( .A1(n648), .A2(n641), .ZN(n645) );
  XOR2_X1 U714 ( .A(KEYINPUT85), .B(KEYINPUT62), .Z(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n646), .A2(n695), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT63), .ZN(G57) );
  INV_X2 U719 ( .A(n648), .ZN(n690) );
  NAND2_X1 U720 ( .A1(n690), .A2(G469), .ZN(n654) );
  XOR2_X1 U721 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n650) );
  XNOR2_X1 U722 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U726 ( .A1(n655), .A2(n695), .ZN(n657) );
  INV_X1 U727 ( .A(KEYINPUT120), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(G54) );
  XNOR2_X1 U729 ( .A(n658), .B(G119), .ZN(G21) );
  NAND2_X1 U730 ( .A1(n690), .A2(G475), .ZN(n662) );
  XOR2_X1 U731 ( .A(KEYINPUT86), .B(KEYINPUT59), .Z(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n663), .A2(n695), .ZN(n665) );
  INV_X1 U735 ( .A(KEYINPUT60), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(G60) );
  XOR2_X1 U737 ( .A(n667), .B(KEYINPUT124), .Z(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n670), .B(n673), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT125), .ZN(n674) );
  XNOR2_X1 U742 ( .A(G227), .B(n674), .ZN(n675) );
  NAND2_X1 U743 ( .A1(G900), .A2(n675), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n676), .A2(G953), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n678), .A2(n677), .ZN(G72) );
  INV_X1 U746 ( .A(n624), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(G953), .ZN(n685) );
  NAND2_X1 U748 ( .A1(G224), .A2(G953), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT123), .ZN(n681) );
  XNOR2_X1 U750 ( .A(n681), .B(KEYINPUT61), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n686), .A2(n687), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n689), .B(n688), .ZN(G69) );
  NAND2_X1 U755 ( .A1(n697), .A2(G217), .ZN(n694) );
  XNOR2_X1 U756 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n691), .B(n692), .ZN(n693) );
  XNOR2_X1 U758 ( .A(n694), .B(n693), .ZN(n696) );
  INV_X1 U759 ( .A(n695), .ZN(n700) );
  NOR2_X1 U760 ( .A1(n696), .A2(n700), .ZN(G66) );
  AND2_X1 U761 ( .A1(n697), .A2(G478), .ZN(n698) );
  XNOR2_X1 U762 ( .A(n699), .B(n698), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n706), .A2(n713), .ZN(n702) );
  XNOR2_X1 U765 ( .A(n702), .B(G104), .ZN(G6) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n704) );
  XNOR2_X1 U767 ( .A(G107), .B(KEYINPUT112), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n704), .B(n703), .ZN(n705) );
  XOR2_X1 U769 ( .A(KEYINPUT26), .B(n705), .Z(n708) );
  NAND2_X1 U770 ( .A1(n706), .A2(n716), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n708), .B(n707), .ZN(G9) );
  XOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .Z(n710) );
  NAND2_X1 U773 ( .A1(n711), .A2(n716), .ZN(n709) );
  XNOR2_X1 U774 ( .A(n710), .B(n709), .ZN(G30) );
  NAND2_X1 U775 ( .A1(n711), .A2(n713), .ZN(n712) );
  XNOR2_X1 U776 ( .A(G146), .B(n712), .ZN(G48) );
  NAND2_X1 U777 ( .A1(n717), .A2(n713), .ZN(n714) );
  XNOR2_X1 U778 ( .A(n714), .B(KEYINPUT114), .ZN(n715) );
  XNOR2_X1 U779 ( .A(G113), .B(n715), .ZN(G15) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U781 ( .A(n718), .B(G116), .ZN(G18) );
  XOR2_X1 U782 ( .A(G125), .B(KEYINPUT37), .Z(n719) );
  XNOR2_X1 U783 ( .A(n720), .B(n719), .ZN(G27) );
  XNOR2_X1 U784 ( .A(G134), .B(n721), .ZN(G36) );
  NAND2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U787 ( .A(KEYINPUT115), .B(n726), .ZN(n728) );
  NAND2_X1 U788 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n748) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n735), .B(KEYINPUT49), .ZN(n736) );
  NAND2_X1 U793 ( .A1(n737), .A2(n736), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n353), .A2(n738), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n740), .B(KEYINPUT50), .ZN(n741) );
  NOR2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U798 ( .A(KEYINPUT51), .B(n745), .Z(n746) );
  NOR2_X1 U799 ( .A1(n752), .A2(n746), .ZN(n747) );
  NOR2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n749), .B(KEYINPUT52), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n754) );
  NOR2_X1 U803 ( .A1(n752), .A2(n731), .ZN(n753) );
  NOR2_X1 U804 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U805 ( .A(KEYINPUT116), .B(n755), .ZN(n762) );
  INV_X1 U806 ( .A(n756), .ZN(n759) );
  NOR2_X1 U807 ( .A1(n757), .A2(KEYINPUT2), .ZN(n758) );
  NOR2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U809 ( .A1(n760), .A2(G953), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U811 ( .A(KEYINPUT117), .B(n763), .ZN(n764) );
  XNOR2_X1 U812 ( .A(KEYINPUT53), .B(n764), .ZN(G75) );
  XOR2_X1 U813 ( .A(n765), .B(G122), .Z(G24) );
  XOR2_X1 U814 ( .A(G137), .B(KEYINPUT126), .Z(n766) );
  XNOR2_X1 U815 ( .A(n767), .B(n766), .ZN(G39) );
  XNOR2_X1 U816 ( .A(G131), .B(KEYINPUT127), .ZN(n769) );
  XNOR2_X1 U817 ( .A(n769), .B(n768), .ZN(G33) );
endmodule

