

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;

  XNOR2_X1 U320 ( .A(n387), .B(KEYINPUT64), .ZN(n388) );
  XNOR2_X1 U321 ( .A(n371), .B(n345), .ZN(n346) );
  XOR2_X1 U322 ( .A(n299), .B(n298), .Z(n580) );
  XOR2_X1 U323 ( .A(n435), .B(KEYINPUT33), .Z(n288) );
  XOR2_X1 U324 ( .A(n293), .B(KEYINPUT31), .Z(n289) );
  XOR2_X1 U325 ( .A(G78GAT), .B(G148GAT), .Z(n290) );
  XNOR2_X1 U326 ( .A(n344), .B(KEYINPUT10), .ZN(n345) );
  INV_X1 U327 ( .A(n351), .ZN(n352) );
  XNOR2_X1 U328 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U329 ( .A(n389), .B(n388), .ZN(n531) );
  XNOR2_X1 U330 ( .A(n355), .B(n354), .ZN(n356) );
  NOR2_X1 U331 ( .A1(n487), .A2(n456), .ZN(n457) );
  NOR2_X1 U332 ( .A1(n534), .A2(n446), .ZN(n572) );
  XNOR2_X1 U333 ( .A(n318), .B(n317), .ZN(n534) );
  XNOR2_X1 U334 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XNOR2_X1 U336 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n290), .B(n291), .ZN(n435) );
  NAND2_X1 U338 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n288), .B(n292), .ZN(n293) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G57GAT), .Z(n419) );
  XNOR2_X1 U341 ( .A(n419), .B(KEYINPUT32), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n289), .B(n294), .ZN(n297) );
  XOR2_X1 U343 ( .A(G64GAT), .B(G92GAT), .Z(n296) );
  XNOR2_X1 U344 ( .A(G176GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n392) );
  XOR2_X1 U346 ( .A(n297), .B(n392), .Z(n299) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .Z(n351) );
  XOR2_X1 U348 ( .A(G71GAT), .B(KEYINPUT13), .Z(n321) );
  XNOR2_X1 U349 ( .A(n351), .B(n321), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n580), .B(KEYINPUT41), .ZN(n379) );
  XOR2_X1 U351 ( .A(n379), .B(KEYINPUT100), .Z(n537) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XOR2_X1 U353 ( .A(G71GAT), .B(KEYINPUT79), .Z(n301) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n303) );
  XOR2_X1 U356 ( .A(G134GAT), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n318) );
  XOR2_X1 U359 ( .A(G176GAT), .B(KEYINPUT20), .Z(n307) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT65), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n316) );
  XOR2_X1 U362 ( .A(G127GAT), .B(KEYINPUT0), .Z(n309) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n406) );
  XOR2_X1 U365 ( .A(G120GAT), .B(n406), .Z(n314) );
  XOR2_X1 U366 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n311) );
  XNOR2_X1 U367 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U369 ( .A(KEYINPUT18), .B(n312), .Z(n399) );
  XNOR2_X1 U370 ( .A(G15GAT), .B(n399), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n317) );
  XOR2_X1 U373 ( .A(G211GAT), .B(G127GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(G8GAT), .B(G183GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n335) );
  XOR2_X1 U376 ( .A(n321), .B(G155GAT), .Z(n324) );
  XNOR2_X1 U377 ( .A(G22GAT), .B(G15GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n322), .B(G1GAT), .ZN(n367) );
  XNOR2_X1 U379 ( .A(n367), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U381 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n326) );
  NAND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U385 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n330) );
  XNOR2_X1 U386 ( .A(KEYINPUT12), .B(G64GAT), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U388 ( .A(G57GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n583) );
  INV_X1 U391 ( .A(n583), .ZN(n560) );
  XOR2_X1 U392 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n337) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n357) );
  XOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  INV_X1 U396 ( .A(G43GAT), .ZN(n338) );
  NAND2_X1 U397 ( .A1(G29GAT), .A2(n338), .ZN(n341) );
  INV_X1 U398 ( .A(G29GAT), .ZN(n339) );
  NAND2_X1 U399 ( .A1(n339), .A2(G43GAT), .ZN(n340) );
  NAND2_X1 U400 ( .A1(n341), .A2(n340), .ZN(n343) );
  XNOR2_X1 U401 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n371) );
  AND2_X1 U403 ( .A1(G232GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U404 ( .A(n397), .B(n346), .Z(n348) );
  XNOR2_X1 U405 ( .A(G92GAT), .B(KEYINPUT66), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n355) );
  XOR2_X1 U407 ( .A(G162GAT), .B(KEYINPUT72), .Z(n350) );
  XNOR2_X1 U408 ( .A(G50GAT), .B(G218GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n439) );
  XOR2_X1 U410 ( .A(G134GAT), .B(KEYINPUT74), .Z(n418) );
  XNOR2_X1 U411 ( .A(n439), .B(n418), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n571) );
  XNOR2_X1 U413 ( .A(n571), .B(KEYINPUT92), .ZN(n359) );
  INV_X1 U414 ( .A(KEYINPUT36), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n487) );
  NOR2_X1 U416 ( .A1(n560), .A2(n487), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(KEYINPUT45), .ZN(n377) );
  XOR2_X1 U418 ( .A(G197GAT), .B(G141GAT), .Z(n362) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G50GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n364) );
  XNOR2_X1 U422 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n375) );
  XOR2_X1 U425 ( .A(G169GAT), .B(G8GAT), .Z(n400) );
  XOR2_X1 U426 ( .A(n367), .B(n400), .Z(n369) );
  NAND2_X1 U427 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U429 ( .A(n370), .B(KEYINPUT29), .Z(n373) );
  XNOR2_X1 U430 ( .A(n371), .B(KEYINPUT68), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n552) );
  INV_X1 U433 ( .A(n552), .ZN(n577) );
  NOR2_X1 U434 ( .A1(n580), .A2(n577), .ZN(n376) );
  AND2_X1 U435 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n378), .B(KEYINPUT107), .ZN(n386) );
  XOR2_X1 U437 ( .A(KEYINPUT106), .B(KEYINPUT47), .Z(n384) );
  NOR2_X1 U438 ( .A1(n379), .A2(n552), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n380), .B(KEYINPUT46), .ZN(n381) );
  NOR2_X1 U440 ( .A1(n583), .A2(n381), .ZN(n382) );
  INV_X1 U441 ( .A(n571), .ZN(n564) );
  NAND2_X1 U442 ( .A1(n382), .A2(n564), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  NAND2_X1 U444 ( .A1(n386), .A2(n385), .ZN(n389) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n387) );
  XOR2_X1 U446 ( .A(KEYINPUT75), .B(KEYINPUT90), .Z(n391) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n396) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(G211GAT), .ZN(n432) );
  XNOR2_X1 U452 ( .A(G218GAT), .B(n432), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U454 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n521) );
  NOR2_X1 U457 ( .A1(n531), .A2(n521), .ZN(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT54), .B(n403), .ZN(n454) );
  XOR2_X1 U459 ( .A(G155GAT), .B(KEYINPUT2), .Z(n405) );
  XNOR2_X1 U460 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n434) );
  XNOR2_X1 U462 ( .A(n406), .B(n434), .ZN(n427) );
  XOR2_X1 U463 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n408) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT85), .B(KEYINPUT88), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U470 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n414) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U473 ( .A(KEYINPUT5), .B(n415), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U475 ( .A(n419), .B(n418), .Z(n421) );
  XNOR2_X1 U476 ( .A(G148GAT), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U478 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G85GAT), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U481 ( .A(n427), .B(n426), .Z(n467) );
  XOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n443) );
  XOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n431) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U488 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U491 ( .A(n438), .B(KEYINPUT81), .Z(n441) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT83), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n469) );
  NOR2_X1 U495 ( .A1(n467), .A2(n469), .ZN(n444) );
  AND2_X1 U496 ( .A1(n454), .A2(n444), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U498 ( .A1(n537), .A2(n572), .ZN(n450) );
  XOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT118), .Z(n448) );
  XNOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n452) );
  XNOR2_X1 U502 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n458) );
  NAND2_X1 U504 ( .A1(n469), .A2(n534), .ZN(n453) );
  XOR2_X1 U505 ( .A(n453), .B(KEYINPUT26), .Z(n550) );
  INV_X1 U506 ( .A(n550), .ZN(n463) );
  INV_X1 U507 ( .A(n467), .ZN(n519) );
  NAND2_X1 U508 ( .A1(n454), .A2(n519), .ZN(n455) );
  NOR2_X2 U509 ( .A1(n463), .A2(n455), .ZN(n584) );
  INV_X1 U510 ( .A(n584), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(n460) );
  INV_X1 U512 ( .A(KEYINPUT124), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(G1355GAT) );
  NOR2_X1 U514 ( .A1(n552), .A2(n580), .ZN(n490) );
  NOR2_X1 U515 ( .A1(n534), .A2(n521), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n469), .A2(n461), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(n462), .Z(n465) );
  XNOR2_X1 U518 ( .A(n521), .B(KEYINPUT27), .ZN(n470) );
  NOR2_X1 U519 ( .A1(n463), .A2(n470), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n474) );
  XOR2_X1 U522 ( .A(KEYINPUT67), .B(KEYINPUT28), .Z(n468) );
  XOR2_X1 U523 ( .A(n469), .B(n468), .Z(n532) );
  INV_X1 U524 ( .A(n532), .ZN(n472) );
  NOR2_X1 U525 ( .A1(n519), .A2(n470), .ZN(n529) );
  NAND2_X1 U526 ( .A1(n529), .A2(n534), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT91), .B(n475), .Z(n486) );
  XOR2_X1 U530 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n477) );
  NAND2_X1 U531 ( .A1(n564), .A2(n583), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n477), .B(n476), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n486), .A2(n478), .ZN(n506) );
  NAND2_X1 U534 ( .A1(n490), .A2(n506), .ZN(n484) );
  NOR2_X1 U535 ( .A1(n519), .A2(n484), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(n479), .Z(n480) );
  XNOR2_X1 U537 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U538 ( .A1(n521), .A2(n484), .ZN(n481) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n534), .A2(n484), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n532), .A2(n484), .ZN(n485) );
  XOR2_X1 U544 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  NOR2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n560), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n489), .ZN(n518) );
  NAND2_X1 U548 ( .A1(n490), .A2(n518), .ZN(n493) );
  XOR2_X1 U549 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n502) );
  NOR2_X1 U552 ( .A1(n519), .A2(n502), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT95), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n496), .Z(G1328GAT) );
  NOR2_X1 U556 ( .A1(n521), .A2(n502), .ZN(n497) );
  XOR2_X1 U557 ( .A(KEYINPUT96), .B(n497), .Z(n498) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n534), .A2(n502), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT97), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U563 ( .A1(n532), .A2(n502), .ZN(n504) );
  XNOR2_X1 U564 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  AND2_X1 U567 ( .A1(n552), .A2(n537), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n517), .A2(n506), .ZN(n512) );
  NOR2_X1 U569 ( .A1(n519), .A2(n512), .ZN(n507) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n512), .ZN(n509) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n534), .A2(n512), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT101), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n532), .ZN(n516) );
  XOR2_X1 U578 ( .A(KEYINPUT103), .B(KEYINPUT43), .Z(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT102), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(n522), .Z(n523) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U588 ( .A1(n534), .A2(n525), .ZN(n524) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT105), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT108), .ZN(n536) );
  INV_X1 U595 ( .A(n529), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n551) );
  NAND2_X1 U597 ( .A1(n551), .A2(n532), .ZN(n533) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n577), .A2(n545), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT49), .B(KEYINPUT109), .Z(n539) );
  NAND2_X1 U602 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n542) );
  NAND2_X1 U607 ( .A1(n545), .A2(n583), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n571), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT112), .Z(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n563) );
  NOR2_X1 U616 ( .A1(n552), .A2(n563), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT114), .B(n554), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n379), .A2(n563), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n556) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT115), .B(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n563), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n577), .A2(n572), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT119), .Z(n568) );
  NAND2_X1 U633 ( .A1(n572), .A2(n583), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT120), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT58), .B(n570), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1351GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT60), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT122), .B(n576), .Z(n579) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT123), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1354GAT) );
endmodule

