//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G77), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n216), .B(new_n217), .C1(new_n203), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G50), .A2(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n202), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT66), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n204), .A2(new_n205), .ZN(new_n233));
  INV_X1    g0033(.A(G50), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n215), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(new_n207), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n231), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n230), .B1(new_n212), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT69), .A2(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT69), .A2(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(new_n231), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n265), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n263), .A2(new_n265), .B1(G50), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(G13), .B(G20), .C1(new_n266), .C2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n234), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(G45), .B1(new_n266), .B2(new_n267), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n268), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G226), .ZN(new_n282));
  INV_X1    g0082(.A(G1), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT68), .B(G45), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(G274), .C1(new_n284), .C2(G41), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G223), .A2(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(new_n276), .C1(G77), .C2(new_n286), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n292), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n297), .B1(new_n298), .B2(new_n292), .C1(new_n275), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n275), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT9), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT10), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT10), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G226), .A2(G1698), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n225), .B2(G1698), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n286), .B1(G33), .B2(G97), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n285), .B1(new_n308), .B2(new_n277), .C1(new_n280), .C2(new_n218), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT13), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(KEYINPUT13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(new_n265), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n272), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n272), .B2(new_n317), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n269), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G68), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n273), .A2(new_n203), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n203), .A2(G20), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n327), .B1(new_n257), .B2(new_n222), .C1(new_n256), .C2(new_n234), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n265), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT74), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n310), .A2(G190), .A3(new_n312), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n316), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n315), .A2(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n315), .A2(new_n339), .A3(G169), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n310), .A2(G179), .A3(new_n312), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n333), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G20), .A2(G77), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT15), .B(G87), .Z(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n345), .B1(new_n260), .B2(new_n256), .C1(new_n257), .C2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n323), .A2(G77), .B1(new_n265), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n273), .A2(new_n222), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G238), .A2(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n286), .B(new_n352), .C1(new_n225), .C2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n276), .C1(G107), .C2(new_n286), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n285), .C1(new_n223), .C2(new_n280), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G200), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n351), .B(new_n356), .C1(new_n298), .C2(new_n355), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n305), .A2(new_n344), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n286), .B2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G33), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n203), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n202), .A2(new_n203), .ZN(new_n368));
  OAI21_X1  g0168(.A(G20), .B1(new_n233), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n255), .A2(G159), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n359), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n359), .C1(new_n367), .C2(new_n371), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n265), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT75), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n363), .A3(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n362), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n360), .A3(new_n231), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n363), .A2(G33), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n377), .B2(new_n379), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT7), .B1(new_n384), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(G68), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n369), .A3(new_n370), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n387), .A2(KEYINPUT76), .A3(new_n359), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT76), .B1(new_n387), .B2(new_n359), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n262), .A2(new_n272), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n270), .B2(new_n262), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n384), .B1(G226), .B2(new_n287), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G223), .A2(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G87), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n395), .A2(new_n396), .B1(new_n264), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n398), .A2(KEYINPUT78), .A3(new_n276), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT78), .B1(new_n398), .B2(new_n276), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n285), .B1(new_n280), .B2(new_n225), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n401), .A2(KEYINPUT79), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(KEYINPUT79), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n399), .A2(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n401), .B1(new_n276), .B2(new_n398), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(G190), .B1(G200), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n394), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n394), .A2(KEYINPUT17), .A3(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n388), .A2(new_n389), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n392), .B1(new_n413), .B2(new_n376), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n404), .A2(G179), .B1(G169), .B2(new_n405), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(KEYINPUT18), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n394), .B2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n351), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n355), .A2(new_n294), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(G179), .C2(new_n355), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n412), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  OR3_X1    g0224(.A1(new_n358), .A2(KEYINPUT80), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT80), .B1(new_n358), .B2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT5), .B(G41), .Z(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n278), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G274), .A3(new_n277), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n384), .A2(G257), .A3(new_n287), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT84), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n365), .A2(G303), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT84), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n384), .A2(new_n436), .A3(G257), .A4(new_n287), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n384), .A2(G264), .A3(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n432), .B1(new_n439), .B2(new_n276), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n430), .A2(new_n276), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G270), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G283), .ZN(new_n444));
  INV_X1    g0244(.A(G97), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n231), .C1(G33), .C2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n265), .C1(new_n231), .C2(G116), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT20), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n273), .ZN(new_n450));
  OAI221_X1 g0250(.A(G116), .B1(new_n264), .B2(new_n268), .C1(new_n319), .C2(new_n321), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n443), .A2(new_n452), .A3(KEYINPUT21), .A4(G169), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n294), .B1(new_n440), .B2(new_n442), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT85), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT21), .A4(new_n452), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n452), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT21), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n443), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n459), .A2(new_n460), .B1(new_n462), .B2(new_n452), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n440), .A2(new_n442), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G190), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n443), .A2(G200), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n450), .A3(new_n451), .A4(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n458), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n384), .B1(G257), .B2(new_n287), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G250), .A2(G1698), .ZN(new_n470));
  INV_X1    g0270(.A(G294), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n469), .A2(new_n470), .B1(new_n264), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n276), .B1(G264), .B2(new_n441), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n431), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G179), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n294), .B2(new_n474), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n384), .A2(KEYINPUT22), .A3(new_n231), .A4(G87), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT86), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(KEYINPUT23), .C1(new_n231), .C2(G107), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n231), .A2(G87), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n365), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT23), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(G20), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT87), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n477), .A2(new_n483), .A3(new_n486), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n265), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n268), .A2(new_n264), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n318), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n272), .A2(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT25), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n476), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n380), .A2(G244), .A3(G1698), .A4(new_n362), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n218), .A2(G1698), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n384), .A2(new_n505), .B1(G33), .B2(G116), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT82), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n384), .A2(new_n507), .A3(G244), .A4(G1698), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n276), .ZN(new_n510));
  INV_X1    g0310(.A(G250), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n278), .B1(KEYINPUT81), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n277), .ZN(new_n513));
  AND2_X1   g0313(.A1(KEYINPUT81), .A2(G250), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n278), .A2(G274), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n510), .A2(new_n461), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n380), .A2(new_n231), .A3(G68), .A4(new_n362), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n520), .A2(new_n264), .A3(new_n445), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G87), .B2(new_n210), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n257), .B2(new_n445), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n519), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n265), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n497), .A2(new_n346), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n273), .A2(new_n347), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n524), .A2(new_n265), .B1(new_n273), .B2(new_n347), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .A3(new_n526), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n518), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n510), .A2(new_n517), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n294), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(G200), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n497), .A2(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n516), .B1(new_n509), .B2(new_n276), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G190), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n533), .A2(new_n535), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n502), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n286), .A2(new_n360), .A3(G20), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT7), .B1(new_n365), .B2(new_n231), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n488), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n445), .A2(new_n488), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n209), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n255), .A2(G77), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n265), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n272), .A2(G97), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n497), .A2(G97), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n286), .B2(G250), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n444), .B(new_n558), .C1(new_n560), .C2(new_n287), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT4), .B1(new_n384), .B2(G244), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n276), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n441), .A2(G257), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n431), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n557), .B(new_n566), .C1(new_n298), .C2(new_n565), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n294), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n563), .A2(new_n461), .A3(new_n431), .A4(new_n564), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n473), .A2(G190), .A3(new_n431), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n495), .A2(new_n573), .A3(new_n498), .A4(new_n500), .ZN(new_n574));
  INV_X1    g0374(.A(G200), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n473), .B2(new_n431), .ZN(new_n576));
  OR3_X1    g0376(.A1(new_n574), .A2(KEYINPUT88), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT88), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n468), .A2(new_n542), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n428), .A2(new_n580), .ZN(G372));
  INV_X1    g0381(.A(new_n296), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n417), .A2(new_n419), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n342), .A2(new_n343), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n336), .B1(new_n584), .B2(new_n423), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n585), .B2(new_n412), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n303), .A2(new_n304), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n582), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT92), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n541), .A2(new_n591), .A3(KEYINPUT26), .A4(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n535), .A2(new_n518), .A3(new_n532), .A4(new_n530), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n539), .A2(G190), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n531), .A2(new_n537), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n536), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n592), .A2(new_n594), .A3(KEYINPUT26), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(KEYINPUT83), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT83), .B1(new_n531), .B2(new_n526), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n510), .A2(KEYINPUT89), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT89), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n509), .A2(new_n605), .A3(new_n276), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n516), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n603), .B(new_n518), .C1(new_n607), .C2(G169), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n540), .B1(new_n607), .B2(new_n575), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n592), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n600), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n518), .A2(new_n530), .A3(new_n532), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n509), .A2(new_n605), .A3(new_n276), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n605), .B1(new_n509), .B2(new_n276), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n517), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n294), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT93), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n595), .A2(new_n596), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(G200), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT90), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n458), .A2(new_n502), .A3(new_n463), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n579), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT91), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n579), .A2(new_n626), .A3(new_n630), .A4(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT93), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT26), .B1(new_n626), .B2(new_n592), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n633), .B(new_n608), .C1(new_n634), .C2(new_n600), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n621), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n590), .B1(new_n428), .B2(new_n637), .ZN(G369));
  NAND2_X1  g0438(.A1(new_n458), .A2(new_n463), .ZN(new_n639));
  INV_X1    g0439(.A(new_n268), .ZN(new_n640));
  INV_X1    g0440(.A(G13), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n639), .A2(new_n452), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT94), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n452), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n468), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(KEYINPUT94), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(G330), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n502), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n501), .A2(new_n648), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT95), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n577), .A2(new_n578), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n502), .A2(new_n648), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n648), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n639), .A2(new_n666), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n662), .A2(new_n667), .B1(new_n502), .B2(new_n648), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n213), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n235), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT98), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n636), .A2(new_n666), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g0482(.A(KEYINPUT98), .B(KEYINPUT29), .C1(new_n636), .C2(new_n666), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n613), .A2(KEYINPUT26), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n608), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n541), .A2(new_n614), .A3(new_n592), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n628), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n666), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT29), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n682), .A2(new_n683), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n468), .A2(new_n542), .A3(new_n579), .A4(new_n666), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n565), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n607), .A2(G179), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n474), .A3(new_n443), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n464), .A2(G179), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n539), .A2(new_n473), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n701), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n462), .A2(KEYINPUT30), .A3(new_n696), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n698), .A2(new_n702), .A3(new_n709), .A4(new_n704), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n648), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n695), .B1(new_n713), .B2(KEYINPUT97), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n666), .B1(new_n705), .B2(KEYINPUT96), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT31), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n717), .B2(new_n707), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n693), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n692), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n678), .B1(new_n720), .B2(G1), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT99), .ZN(G364));
  NAND2_X1  g0522(.A1(new_n642), .A2(G45), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n673), .A2(G1), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n654), .A2(G20), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n230), .B1(G20), .B2(new_n294), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(G355), .A2(new_n286), .A3(new_n213), .ZN(new_n731));
  INV_X1    g0531(.A(G45), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n248), .A2(new_n732), .B1(new_n676), .B2(new_n284), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n384), .A2(new_n671), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n731), .B1(G116), .B2(new_n213), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n724), .B(new_n727), .C1(new_n730), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n461), .A2(new_n575), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n231), .A2(new_n298), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n234), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n575), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n397), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n231), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G159), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT32), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n461), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n745), .A2(new_n742), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n222), .A2(new_n752), .B1(new_n753), .B2(new_n488), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n231), .B1(new_n746), .B2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n739), .A2(new_n751), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n286), .B1(new_n755), .B2(new_n445), .C1(new_n202), .C2(new_n756), .ZN(new_n757));
  OR4_X1    g0557(.A1(new_n744), .A2(new_n750), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n738), .A2(new_n745), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n741), .B(new_n758), .C1(G68), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G317), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(KEYINPUT33), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n748), .A2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n753), .ZN(new_n768));
  INV_X1    g0568(.A(new_n740), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(G326), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n743), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G303), .ZN(new_n772));
  INV_X1    g0572(.A(new_n756), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n286), .B1(new_n773), .B2(G322), .ZN(new_n774));
  INV_X1    g0574(.A(new_n755), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G294), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n770), .A2(new_n772), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n752), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(G311), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n729), .B1(new_n761), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n654), .A2(G330), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n724), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n656), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n737), .A2(new_n780), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  OR2_X1    g0586(.A1(new_n423), .A2(new_n648), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n357), .B1(new_n351), .B2(new_n666), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n423), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n636), .A2(new_n666), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n636), .B2(new_n666), .ZN(new_n795));
  OR3_X1    g0595(.A1(new_n794), .A2(new_n719), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n719), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(new_n724), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n729), .A2(new_n725), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n222), .ZN(new_n800));
  INV_X1    g0600(.A(G137), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n740), .A2(new_n801), .B1(new_n759), .B2(new_n254), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT101), .Z(new_n803));
  AOI22_X1  g0603(.A1(G143), .A2(new_n773), .B1(new_n778), .B2(G159), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT34), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(KEYINPUT34), .A3(new_n804), .ZN(new_n806));
  INV_X1    g0606(.A(new_n753), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G68), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n743), .A2(new_n234), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n381), .B(new_n809), .C1(G132), .C2(new_n748), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n805), .B(new_n811), .C1(G58), .C2(new_n775), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n807), .A2(G87), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n471), .B2(new_n756), .C1(new_n814), .C2(new_n747), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G107), .B2(new_n771), .ZN(new_n816));
  INV_X1    g0616(.A(G303), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n740), .A2(new_n817), .B1(new_n755), .B2(new_n445), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n286), .B(new_n818), .C1(G116), .C2(new_n778), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n816), .B(new_n819), .C1(new_n767), .C2(new_n759), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT100), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n729), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n800), .B(new_n822), .C1(new_n792), .C2(new_n726), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n798), .B1(new_n724), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT102), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G384));
  NAND2_X1  g0627(.A1(new_n388), .A2(new_n389), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n317), .B1(new_n387), .B2(new_n359), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n392), .ZN(new_n831));
  INV_X1    g0631(.A(new_n646), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n407), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n415), .B1(new_n830), .B2(new_n392), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT104), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n414), .A2(new_n837), .A3(new_n416), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT104), .B1(new_n394), .B2(new_n415), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n414), .A2(new_n832), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n407), .ZN(new_n841));
  XOR2_X1   g0641(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n842));
  OAI21_X1  g0642(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n832), .B(new_n831), .C1(new_n583), .C2(new_n411), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n840), .A2(new_n407), .ZN(new_n846));
  INV_X1    g0646(.A(new_n842), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(new_n838), .A4(new_n839), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n840), .A2(new_n407), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n394), .A2(new_n415), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n420), .A2(new_n409), .A3(new_n410), .ZN(new_n852));
  INV_X1    g0652(.A(new_n840), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n848), .A2(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n845), .B1(new_n854), .B2(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n343), .A2(new_n648), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n344), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n584), .B2(new_n666), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n711), .A2(new_n712), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n694), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n855), .A2(new_n792), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AND4_X1   g0663(.A1(new_n863), .A2(new_n858), .A3(new_n861), .A4(new_n792), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n843), .A2(new_n844), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n845), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n862), .A2(KEYINPUT40), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n427), .A2(new_n861), .ZN(new_n871));
  OAI21_X1  g0671(.A(G330), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n680), .A2(new_n681), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT98), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n680), .A2(new_n679), .A3(new_n681), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(new_n427), .A3(new_n690), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n682), .A2(new_n683), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT107), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n427), .A4(new_n690), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n589), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n873), .B(new_n882), .Z(new_n883));
  INV_X1    g0683(.A(KEYINPUT106), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n848), .A2(new_n851), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n852), .A2(new_n853), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n887), .B2(new_n866), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n868), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n866), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(new_n884), .A3(new_n891), .A4(new_n845), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n584), .A2(new_n648), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n893), .A2(new_n894), .B1(new_n583), .B2(new_n646), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n793), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n868), .A3(new_n858), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n883), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n640), .B2(new_n642), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n449), .B1(new_n549), .B2(KEYINPUT35), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n232), .C1(KEYINPUT35), .C2(new_n549), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  OAI21_X1  g0705(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n676), .A2(new_n906), .B1(G50), .B2(new_n203), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n641), .A3(new_n268), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NOR2_X1   g0709(.A1(new_n666), .A2(new_n596), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n608), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n626), .B2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n728), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n753), .A2(new_n445), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n743), .A2(new_n449), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT46), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT116), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n769), .A2(G311), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n752), .A2(new_n767), .B1(new_n755), .B2(new_n488), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT115), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n759), .A2(new_n471), .B1(new_n747), .B2(new_n762), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n384), .B(new_n922), .C1(KEYINPUT46), .C2(new_n916), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n918), .A2(new_n919), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n915), .B(new_n924), .C1(G303), .C2(new_n773), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n778), .A2(G50), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n769), .A2(G143), .B1(new_n775), .B2(G68), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n254), .B2(new_n756), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n928), .A2(KEYINPUT117), .B1(new_n222), .B2(new_n753), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT117), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n743), .A2(new_n202), .B1(new_n747), .B2(new_n801), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n365), .B1(new_n931), .B2(KEYINPUT118), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n930), .B(new_n932), .C1(KEYINPUT118), .C2(new_n931), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n929), .B(new_n933), .C1(G159), .C2(new_n760), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n925), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT47), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n729), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n730), .B1(new_n213), .B2(new_n347), .C1(new_n239), .C2(new_n735), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n914), .A2(new_n783), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n723), .A2(G1), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT114), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n557), .A2(new_n666), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n572), .A2(new_n942), .B1(new_n571), .B2(new_n666), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT109), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n668), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT44), .Z(new_n947));
  INV_X1    g0747(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT112), .B1(new_n668), .B2(new_n945), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n668), .A2(new_n945), .A3(KEYINPUT112), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n947), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT113), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n665), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT113), .B1(new_n958), .B2(KEYINPUT114), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n957), .A2(new_n958), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n667), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n664), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n655), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n720), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n672), .B(KEYINPUT41), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n940), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n913), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n592), .B1(new_n944), .B2(new_n657), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT110), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n666), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n664), .A2(new_n961), .A3(new_n944), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT42), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n968), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n913), .A2(new_n967), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT111), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n665), .B2(new_n945), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n665), .A2(new_n945), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n939), .B1(new_n966), .B2(new_n983), .ZN(G387));
  INV_X1    g0784(.A(new_n963), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n720), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n963), .B1(new_n692), .B2(new_n719), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n672), .A3(new_n987), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n260), .A2(KEYINPUT50), .A3(G50), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT50), .B1(new_n260), .B2(G50), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(new_n732), .A4(new_n674), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G68), .B2(G77), .ZN(new_n992));
  INV_X1    g0792(.A(new_n284), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n734), .B1(new_n243), .B2(new_n993), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n674), .A2(new_n671), .A3(new_n365), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n213), .A2(G107), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n998), .A2(new_n729), .A3(new_n728), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n664), .A2(G20), .A3(new_n726), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G50), .A2(new_n773), .B1(new_n748), .B2(G150), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n347), .B2(new_n755), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n915), .B(new_n1002), .C1(G159), .C2(new_n769), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n771), .A2(G77), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n778), .A2(G68), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n381), .B1(new_n261), .B2(new_n760), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n771), .A2(G294), .B1(new_n775), .B2(G283), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n756), .A2(new_n762), .B1(new_n752), .B2(new_n817), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT119), .ZN(new_n1010));
  INV_X1    g0810(.A(G322), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n814), .B2(new_n759), .C1(new_n1011), .C2(new_n740), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT48), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1008), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT120), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n748), .A2(G326), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n807), .A2(G116), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1017), .A2(new_n381), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1007), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n999), .B(new_n1000), .C1(new_n1022), .C2(new_n729), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n985), .A2(new_n940), .B1(new_n1023), .B2(new_n783), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n988), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT121), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n988), .A2(KEYINPUT121), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(G393));
  AND2_X1   g0829(.A1(new_n954), .A2(new_n952), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT122), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n958), .A4(new_n947), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n958), .A2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n665), .A2(KEYINPUT122), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n955), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n986), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n672), .C1(new_n960), .C2(new_n986), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n740), .A2(new_n762), .B1(new_n756), .B2(new_n814), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT52), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n365), .B1(new_n753), .B2(new_n488), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n759), .A2(new_n817), .B1(new_n747), .B2(new_n1011), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n743), .A2(new_n767), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n449), .B2(new_n755), .C1(new_n471), .C2(new_n752), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT124), .Z(new_n1045));
  NOR2_X1   g0845(.A1(new_n752), .A2(new_n260), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n759), .A2(new_n234), .B1(new_n755), .B2(new_n222), .ZN(new_n1047));
  INV_X1    g0847(.A(G159), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n740), .A2(new_n254), .B1(new_n756), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT51), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n1047), .B(new_n1050), .C1(G68), .C2(new_n771), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n381), .B1(G143), .B2(new_n748), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n813), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT125), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n729), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n730), .B1(new_n445), .B2(new_n213), .C1(new_n251), .C2(new_n735), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n724), .B1(new_n945), .B2(new_n728), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1032), .A2(KEYINPUT123), .A3(new_n1035), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT123), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n940), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1037), .A2(new_n1059), .A3(new_n1063), .ZN(G390));
  AND2_X1   g0864(.A1(new_n889), .A2(new_n892), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n725), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n752), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n759), .A2(new_n801), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n365), .B(new_n1069), .C1(G132), .C2(new_n773), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n775), .A2(G159), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n743), .A2(new_n254), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT53), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G50), .A2(new_n807), .B1(new_n748), .B2(G125), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1068), .B(new_n1075), .C1(G128), .C2(new_n769), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n752), .A2(new_n445), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n744), .B1(G68), .B2(new_n807), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n769), .A2(G283), .B1(new_n748), .B2(G294), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n286), .B1(new_n775), .B2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n760), .A2(G107), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1077), .B(new_n1082), .C1(G116), .C2(new_n773), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n729), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1066), .A2(new_n783), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n262), .B2(new_n799), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n718), .A3(new_n694), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1088), .A2(G330), .A3(new_n792), .A4(new_n858), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT126), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT126), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n719), .A2(new_n1091), .A3(new_n792), .A4(new_n858), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n894), .B1(new_n890), .B2(new_n845), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n787), .B1(new_n688), .B2(new_n791), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n858), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n894), .B1(new_n898), .B2(new_n858), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1093), .B(new_n1097), .C1(new_n893), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n898), .A2(new_n858), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n894), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(new_n1065), .B1(new_n1096), .B2(new_n1094), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n861), .A2(new_n792), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n858), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n693), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1099), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1086), .B1(new_n1109), .B2(new_n940), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n427), .A2(G330), .A3(new_n861), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1095), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1105), .B1(new_n1104), .B2(new_n693), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1093), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n858), .B1(new_n719), .B2(new_n792), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n898), .B1(new_n1116), .B2(new_n1106), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n882), .A2(new_n1112), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n1109), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n672), .B1(new_n1119), .B2(new_n1108), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(G378));
  XOR2_X1   g0923(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n305), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n305), .A2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n301), .A2(new_n646), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n725), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n753), .A2(new_n202), .B1(new_n747), .B2(new_n767), .ZN(new_n1134));
  AOI21_X1  g0934(.A(G41), .B1(new_n769), .B2(G116), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n778), .A2(new_n346), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1135), .A2(new_n381), .A3(new_n1004), .A4(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1134), .B(new_n1137), .C1(G68), .C2(new_n775), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n445), .B2(new_n759), .C1(new_n488), .C2(new_n756), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT58), .Z(new_n1140));
  OAI22_X1  g0940(.A1(new_n743), .A2(new_n1067), .B1(new_n755), .B2(new_n254), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n756), .A2(new_n1142), .B1(new_n752), .B2(new_n801), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(G125), .C2(new_n769), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n760), .A2(G132), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT59), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G33), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n748), .B2(G124), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n1048), .C2(new_n753), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G41), .B1(new_n380), .B2(G33), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1150), .A2(new_n1151), .B1(G50), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n729), .B1(new_n1140), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n799), .A2(new_n234), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n783), .A2(new_n1133), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n869), .B2(new_n693), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n864), .A2(new_n868), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n863), .B1(new_n1160), .B2(new_n855), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n1132), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  AND4_X1   g0962(.A1(new_n899), .A2(new_n1158), .A3(new_n895), .A4(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1158), .A2(new_n1162), .B1(new_n895), .B2(new_n899), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1165), .B2(new_n940), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n589), .B(new_n1111), .C1(new_n878), .C2(new_n881), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1108), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(KEYINPUT57), .A3(new_n1165), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n672), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1165), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(G375));
  AOI21_X1  g0973(.A(new_n1118), .B1(new_n882), .B2(new_n1112), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n965), .A3(new_n1119), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n759), .A2(new_n449), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G77), .A2(new_n807), .B1(new_n778), .B2(G107), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n769), .A2(G294), .B1(new_n775), .B2(new_n346), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n748), .A2(G303), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n286), .B1(new_n771), .B2(G97), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1177), .B(new_n1182), .C1(G283), .C2(new_n773), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G132), .A2(new_n769), .B1(new_n771), .B2(G159), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n234), .B2(new_n755), .C1(new_n254), .C2(new_n752), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n747), .A2(new_n1142), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n759), .A2(new_n1067), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n384), .B1(new_n753), .B2(new_n202), .C1(new_n801), .C2(new_n756), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n729), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n783), .B(new_n1190), .C1(new_n858), .C2(new_n726), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n203), .B2(new_n799), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1118), .B2(new_n940), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1176), .A2(new_n1193), .ZN(G381));
  OR2_X1    g0994(.A1(G375), .A2(G378), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1195), .A2(G384), .A3(G381), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G387), .A2(G390), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1027), .A2(new_n785), .A3(new_n1028), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(G407));
  INV_X1    g1000(.A(G213), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(G343), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1195), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(KEYINPUT127), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G407), .B(new_n1205), .C1(KEYINPUT127), .C2(new_n1204), .ZN(G409));
  NAND2_X1  g1006(.A1(G375), .A2(G378), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n672), .B(new_n1119), .C1(new_n1174), .C2(KEYINPUT60), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n878), .A2(new_n881), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n590), .A3(new_n1112), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(KEYINPUT60), .A3(new_n1168), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1193), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G384), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1167), .B2(new_n1118), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(new_n672), .A3(new_n1211), .A4(new_n1119), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n826), .A3(new_n1193), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1169), .A2(new_n965), .A3(new_n1165), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1166), .ZN(new_n1221));
  OR2_X1    g1021(.A1(G378), .A2(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1207), .A2(new_n1219), .A3(new_n1203), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1202), .B1(G375), .B2(G378), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1202), .A2(G2897), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1217), .A2(new_n826), .A3(new_n1193), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n826), .B1(new_n1217), .B2(new_n1193), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1214), .A2(new_n1218), .A3(new_n1225), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1224), .A2(new_n1222), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT63), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1223), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  AND2_X1   g1034(.A1(G387), .A2(G390), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1198), .B(new_n1234), .C1(new_n1235), .C2(new_n1197), .ZN(new_n1236));
  OR2_X1    g1036(.A1(G387), .A2(G390), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1198), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(G390), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1224), .A2(KEYINPUT63), .A3(new_n1219), .A4(new_n1222), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1223), .A2(KEYINPUT62), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1207), .A2(new_n1203), .A3(new_n1222), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1223), .B2(KEYINPUT62), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1246), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1245), .A2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(new_n1195), .A2(new_n1207), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1241), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1246), .A2(new_n1195), .A3(new_n1207), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1219), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1218), .A3(new_n1257), .A4(new_n1214), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(G402));
endmodule


