//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(new_n467), .A3(G101), .A4(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n466), .A2(G137), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n464), .B2(new_n465), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n467), .B1(new_n464), .B2(new_n465), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n481), .B(new_n483), .C1(G124), .C2(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n484), .A2(G126), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n467), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n495), .A2(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n506), .B(KEYINPUT71), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n503), .B2(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n503), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G88), .B1(new_n517), .B2(G50), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n512), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n511), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n522), .A2(new_n503), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n530), .A2(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR3_X1    g112(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n533), .B2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n515), .A2(G81), .B1(new_n517), .B2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT73), .Z(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n517), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n531), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n503), .B(KEYINPUT74), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G65), .Z(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(new_n556), .B1(G78), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  OR3_X1    g133(.A1(new_n557), .A2(new_n558), .A3(new_n536), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n557), .B2(new_n536), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n515), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n517), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n536), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n515), .A2(G86), .B1(new_n517), .B2(G48), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G305));
  AND2_X1   g150(.A1(new_n503), .A2(G60), .ZN(new_n576));
  AND2_X1   g151(.A1(G72), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n515), .A2(G85), .B1(new_n517), .B2(G47), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G301), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n515), .A2(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G54), .B2(new_n517), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n555), .A2(G66), .ZN(new_n589));
  AND2_X1   g164(.A1(G79), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(new_n584), .ZN(G284));
  XOR2_X1   g169(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n561), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(new_n561), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n593), .B1(new_n599), .B2(G860), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n545), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g181(.A1(new_n467), .A2(G2104), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n493), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n466), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n484), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n467), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n631), .ZN(G401));
  XOR2_X1   g211(.A(G2067), .B(G2678), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT84), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n639), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n639), .B(KEYINPUT17), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n644), .B(new_n641), .C1(new_n638), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n638), .A3(new_n640), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  AOI211_X1 g234(.A(new_n657), .B(new_n659), .C1(new_n652), .C2(new_n656), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1981), .B(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G229));
  INV_X1    g241(.A(G16), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G23), .ZN(new_n668));
  XNOR2_X1  g243(.A(G288), .B(KEYINPUT86), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n669), .B2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT33), .Z(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(G1976), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(G1976), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(G22), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G166), .B2(new_n667), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1971), .ZN(new_n676));
  MUX2_X1   g251(.A(G6), .B(G305), .S(G16), .Z(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  NOR4_X1   g254(.A1(new_n672), .A2(new_n673), .A3(new_n676), .A4(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n684));
  INV_X1    g259(.A(G107), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G2105), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  AOI22_X1  g262(.A1(G119), .A2(new_n484), .B1(new_n466), .B2(G131), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  MUX2_X1   g264(.A(G25), .B(new_n689), .S(G29), .Z(new_n690));
  XOR2_X1   g265(.A(KEYINPUT35), .B(G1991), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n667), .A2(G24), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G290), .B2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n682), .A2(new_n683), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT36), .ZN(new_n699));
  NOR2_X1   g274(.A1(G4), .A2(G16), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n593), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G2090), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G35), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n703), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT29), .Z(new_n707));
  AOI22_X1  g282(.A1(new_n701), .A2(G1348), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G5), .A2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G171), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT89), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n703), .A2(G32), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n466), .A2(G141), .B1(G105), .B2(new_n607), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n484), .A2(G129), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT26), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n703), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n708), .B1(G1961), .B2(new_n711), .C1(new_n713), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n713), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT90), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n667), .A2(G20), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n561), .B2(new_n667), .ZN(new_n729));
  INV_X1    g304(.A(G1956), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n667), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n545), .B2(new_n667), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1341), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n701), .A2(G1348), .B1(new_n702), .B2(new_n707), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n711), .A2(G1961), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n703), .A2(G27), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT93), .Z(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n703), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(KEYINPUT24), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n477), .B2(new_n703), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n739), .A2(G2078), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n703), .A2(G33), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n747));
  NAND2_X1  g322(.A1(G103), .A2(G2104), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2105), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n466), .A2(G139), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n467), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n736), .B(new_n745), .C1(new_n442), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n739), .A2(G2078), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n754), .A2(new_n442), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT91), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n703), .B1(new_n760), .B2(G28), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n759), .B1(new_n761), .B2(new_n762), .C1(new_n618), .C2(new_n703), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n744), .A2(new_n740), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n756), .A2(new_n757), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n703), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G116), .B2(new_n467), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT87), .ZN(new_n771));
  AOI22_X1  g346(.A1(G128), .A2(new_n484), .B1(new_n466), .B2(G140), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n703), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n667), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n667), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n765), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n734), .A2(new_n735), .A3(new_n755), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n726), .A2(new_n731), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT95), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n699), .A2(new_n784), .ZN(G150));
  INV_X1    g360(.A(G150), .ZN(G311));
  NAND2_X1  g361(.A1(new_n515), .A2(G93), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT96), .B(G55), .Z(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n536), .B2(new_n788), .C1(new_n523), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n543), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT38), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n593), .A2(G559), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT39), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(KEYINPUT39), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n797), .A2(new_n798), .A3(G860), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n790), .A2(G860), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT37), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n801), .ZN(G145));
  INV_X1    g377(.A(KEYINPUT103), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n484), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n487), .B1(new_n490), .B2(new_n489), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT4), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n806), .A2(KEYINPUT99), .A3(new_n491), .ZN(new_n807));
  AOI21_X1  g382(.A(KEYINPUT99), .B1(new_n806), .B2(new_n491), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(KEYINPUT100), .B(new_n804), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n773), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(new_n719), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n719), .ZN(new_n817));
  OAI211_X1 g392(.A(KEYINPUT101), .B(new_n753), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n753), .A2(KEYINPUT101), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n753), .A2(KEYINPUT101), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n815), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n689), .B(new_n609), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n466), .A2(G142), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n484), .A2(G130), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n467), .A2(G118), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n824), .B(new_n829), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n830), .B1(new_n818), .B2(new_n822), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(G162), .B(new_n477), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n618), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(G37), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n823), .B(new_n831), .ZN(new_n841));
  INV_X1    g416(.A(new_n838), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n842), .C1(new_n832), .C2(new_n833), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n803), .B(new_n839), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n842), .B1(new_n832), .B2(new_n833), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT102), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n844), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n803), .B1(new_n850), .B2(new_n839), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n847), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n839), .B1(new_n843), .B2(new_n845), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT103), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT40), .B1(new_n855), .B2(new_n846), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(G395));
  NAND2_X1  g432(.A1(new_n790), .A2(new_n584), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n602), .B(KEYINPUT104), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n793), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n593), .A2(G299), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n592), .A2(new_n561), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n593), .A2(KEYINPUT105), .A3(G299), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(KEYINPUT41), .A3(new_n865), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n861), .A2(new_n869), .A3(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n860), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT106), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n669), .B(G303), .ZN(new_n873));
  XOR2_X1   g448(.A(G290), .B(G305), .Z(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT42), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n867), .A2(KEYINPUT106), .A3(new_n871), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n858), .B1(new_n879), .B2(new_n584), .ZN(G295));
  OAI21_X1  g455(.A(new_n858), .B1(new_n879), .B2(new_n584), .ZN(G331));
  NAND2_X1  g456(.A1(new_n868), .A2(new_n870), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n883));
  AOI21_X1  g458(.A(G286), .B1(G171), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(G171), .A2(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n886), .B2(new_n887), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n891), .A2(new_n892), .A3(new_n793), .ZN(new_n893));
  INV_X1    g468(.A(new_n793), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n887), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n888), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n896), .B2(new_n890), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n882), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n793), .B1(new_n891), .B2(new_n892), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n890), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(new_n866), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n875), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n875), .A3(new_n901), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT109), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n910), .A3(KEYINPUT43), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n869), .B1(new_n899), .B2(new_n900), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n861), .A2(new_n863), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n866), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n912), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n902), .B2(new_n903), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n909), .A2(new_n911), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n907), .A2(new_n918), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  MUX2_X1   g498(.A(new_n920), .B(new_n923), .S(KEYINPUT44), .Z(G397));
  NAND3_X1  g499(.A1(new_n472), .A2(new_n476), .A3(G40), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT110), .Z(new_n926));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT45), .B(new_n926), .C1(new_n813), .C2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n773), .B(G2067), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n719), .B(G1996), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n687), .A2(new_n691), .A3(new_n688), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G290), .B(G1986), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n928), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G8), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n925), .B(KEYINPUT110), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n927), .B1(new_n495), .B2(new_n501), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT50), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n809), .A2(new_n927), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n940), .B(new_n942), .C1(new_n943), .C2(KEYINPUT50), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n740), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n806), .A2(new_n491), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n947), .B2(new_n804), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n949));
  INV_X1    g524(.A(new_n943), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n940), .B(new_n949), .C1(new_n950), .C2(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n779), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n939), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT51), .B1(new_n953), .B2(KEYINPUT124), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n946), .A2(G168), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G8), .ZN(new_n957));
  AOI21_X1  g532(.A(G168), .B1(new_n946), .B2(new_n952), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT62), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n959), .B(new_n960), .C1(new_n955), .C2(new_n957), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n955), .A2(new_n957), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n957), .A2(new_n958), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n954), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT62), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n945), .A2(G1961), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n811), .A2(new_n812), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n812), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n941), .B2(new_n968), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n948), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n940), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n967), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT113), .B(new_n978), .C1(new_n972), .C2(new_n973), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n443), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n966), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n951), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n961), .A2(new_n965), .A3(G171), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n972), .B2(new_n973), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(new_n442), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n561), .B(KEYINPUT57), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n948), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT118), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n995), .B(new_n940), .C1(new_n993), .C2(new_n950), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n730), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n926), .A2(new_n943), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n775), .ZN(new_n1001));
  INV_X1    g576(.A(G1348), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n944), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n593), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT122), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n991), .A2(new_n997), .ZN(new_n1007));
  INV_X1    g582(.A(new_n992), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n999), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n998), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n974), .A2(new_n979), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT58), .B(G1341), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1000), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n545), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT123), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n1004), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1001), .A2(new_n1003), .A3(KEYINPUT123), .A4(KEYINPUT60), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n592), .B1(new_n1004), .B2(new_n1021), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT59), .B(new_n545), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1025), .A3(new_n1023), .ZN(new_n1029));
  AND4_X1   g604(.A1(new_n1019), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1010), .B1(new_n1012), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(G171), .B(KEYINPUT54), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n986), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n959), .B1(new_n955), .B2(new_n957), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n813), .B2(new_n927), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(new_n925), .A3(new_n985), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1036), .B2(new_n974), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n984), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n987), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n669), .A2(G1976), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(G8), .C1(new_n926), .C2(new_n943), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(new_n1043), .B2(KEYINPUT116), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(KEYINPUT116), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1000), .A2(new_n939), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1049));
  OR2_X1    g624(.A1(G305), .A2(G1981), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n571), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1046), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1045), .A2(new_n1049), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1061));
  INV_X1    g636(.A(G1971), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n988), .A2(new_n967), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(G2090), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n944), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n939), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G166), .A2(new_n939), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1070), .B(KEYINPUT55), .Z(new_n1071));
  XOR2_X1   g646(.A(new_n1071), .B(KEYINPUT115), .Z(new_n1072));
  AOI21_X1  g647(.A(new_n1060), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n996), .A2(new_n1066), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n980), .A2(new_n981), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1062), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1076), .B2(new_n939), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1040), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G288), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1059), .A2(new_n1047), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1050), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1046), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G8), .A3(new_n1072), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1085), .B2(new_n1060), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1060), .ZN(new_n1087));
  INV_X1    g662(.A(new_n953), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(G286), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1077), .A2(new_n1085), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1073), .A2(KEYINPUT119), .A3(new_n1077), .A4(new_n1089), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1088), .A2(new_n1093), .A3(G286), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1071), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1073), .B(new_n1096), .C1(new_n1097), .C2(new_n1069), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1086), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1079), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT120), .B(new_n1086), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n938), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1996), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n928), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT46), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n928), .B1(new_n719), .B2(new_n930), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT47), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n936), .A2(new_n928), .ZN(new_n1112));
  NOR2_X1   g687(.A1(G290), .A2(G1986), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n928), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT48), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1115), .B2(new_n1114), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n773), .A2(new_n775), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n934), .B(KEYINPUT125), .Z(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n933), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n928), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1111), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1103), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g701(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1128));
  OAI211_X1 g702(.A(new_n920), .B(new_n1128), .C1(new_n847), .C2(new_n851), .ZN(G225));
  INV_X1    g703(.A(G225), .ZN(G308));
endmodule


