

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X1 U324 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U325 ( .A(n311), .B(n310), .Z(n568) );
  XOR2_X1 U326 ( .A(KEYINPUT45), .B(n371), .Z(n292) );
  XNOR2_X1 U327 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n401) );
  XNOR2_X1 U328 ( .A(n402), .B(n401), .ZN(n403) );
  INV_X1 U329 ( .A(KEYINPUT64), .ZN(n445) );
  XNOR2_X1 U330 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U331 ( .A(KEYINPUT77), .B(G64GAT), .Z(n417) );
  XOR2_X1 U332 ( .A(KEYINPUT84), .B(n568), .Z(n486) );
  XOR2_X1 U333 ( .A(n464), .B(n463), .Z(n531) );
  XNOR2_X1 U334 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U335 ( .A(n469), .B(n468), .ZN(G1351GAT) );
  XNOR2_X1 U336 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n293), .B(KEYINPUT83), .ZN(n420) );
  XOR2_X1 U338 ( .A(n420), .B(KEYINPUT82), .Z(n295) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n311) );
  XOR2_X1 U341 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n297) );
  XNOR2_X1 U342 ( .A(KEYINPUT81), .B(KEYINPUT66), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n298), .B(KEYINPUT80), .Z(n300) );
  XOR2_X1 U345 ( .A(G43GAT), .B(G134GAT), .Z(n451) );
  XNOR2_X1 U346 ( .A(n451), .B(KEYINPUT10), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U348 ( .A(KEYINPUT76), .B(G92GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(G106GAT), .B(n303), .Z(n390) );
  XNOR2_X1 U352 ( .A(n304), .B(n390), .ZN(n309) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n305), .B(KEYINPUT8), .ZN(n343) );
  XOR2_X1 U355 ( .A(G162GAT), .B(KEYINPUT79), .Z(n307) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n324) );
  XOR2_X1 U358 ( .A(n343), .B(n324), .Z(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U360 ( .A(G211GAT), .B(KEYINPUT97), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n312), .B(KEYINPUT21), .ZN(n313) );
  XOR2_X1 U362 ( .A(n313), .B(KEYINPUT96), .Z(n315) );
  XNOR2_X1 U363 ( .A(G197GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n414) );
  XOR2_X1 U365 ( .A(G22GAT), .B(G155GAT), .Z(n360) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n316), .B(KEYINPUT2), .ZN(n431) );
  XOR2_X1 U368 ( .A(n360), .B(n431), .Z(n318) );
  XNOR2_X1 U369 ( .A(G106GAT), .B(KEYINPUT22), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n414), .B(n319), .ZN(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT98), .B(KEYINPUT23), .Z(n321) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n322), .B(KEYINPUT24), .Z(n326) );
  XNOR2_X1 U376 ( .A(G78GAT), .B(KEYINPUT75), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n323), .B(G148GAT), .ZN(n391) );
  XNOR2_X1 U378 ( .A(n324), .B(n391), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n480) );
  XOR2_X1 U381 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n330) );
  XNOR2_X1 U382 ( .A(G15GAT), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n342) );
  XOR2_X1 U384 ( .A(G197GAT), .B(G50GAT), .Z(n332) );
  XNOR2_X1 U385 ( .A(G43GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n340) );
  XOR2_X1 U387 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n334) );
  XNOR2_X1 U388 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G22GAT), .Z(n336) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G141GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U393 ( .A(n338), .B(n337), .Z(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U396 ( .A(G1GAT), .B(KEYINPUT70), .Z(n361) );
  XOR2_X1 U397 ( .A(n343), .B(n361), .Z(n345) );
  NAND2_X1 U398 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U400 ( .A(n347), .B(n346), .Z(n559) );
  INV_X1 U401 ( .A(n559), .ZN(n582) );
  XOR2_X1 U402 ( .A(KEYINPUT86), .B(KEYINPUT14), .Z(n349) );
  XNOR2_X1 U403 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n369) );
  XOR2_X1 U405 ( .A(G78GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U406 ( .A(G183GAT), .B(G71GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U408 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n353) );
  XNOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT89), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U411 ( .A(n355), .B(n354), .Z(n367) );
  XOR2_X1 U412 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n357) );
  XNOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n387) );
  XOR2_X1 U415 ( .A(n387), .B(KEYINPUT87), .Z(n359) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U418 ( .A(G8GAT), .B(KEYINPUT85), .Z(n419) );
  XOR2_X1 U419 ( .A(n419), .B(n360), .Z(n363) );
  XOR2_X1 U420 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XNOR2_X1 U421 ( .A(n361), .B(n449), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n590) );
  INV_X1 U426 ( .A(n590), .ZN(n577) );
  XOR2_X1 U427 ( .A(KEYINPUT36), .B(KEYINPUT105), .Z(n370) );
  XNOR2_X1 U428 ( .A(n486), .B(n370), .ZN(n593) );
  NOR2_X1 U429 ( .A1(n577), .A2(n593), .ZN(n371) );
  INV_X1 U430 ( .A(n417), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n372), .A2(G204GAT), .ZN(n375) );
  INV_X1 U432 ( .A(G204GAT), .ZN(n373) );
  NAND2_X1 U433 ( .A1(n417), .A2(n373), .ZN(n374) );
  NAND2_X1 U434 ( .A1(n375), .A2(n374), .ZN(n377) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(n450), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n383) );
  INV_X1 U438 ( .A(n383), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n378) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n382) );
  INV_X1 U442 ( .A(n382), .ZN(n380) );
  NAND2_X1 U443 ( .A1(n381), .A2(n380), .ZN(n385) );
  NAND2_X1 U444 ( .A1(n383), .A2(n382), .ZN(n384) );
  NAND2_X1 U445 ( .A1(n385), .A2(n384), .ZN(n389) );
  AND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n395) );
  NOR2_X1 U449 ( .A1(n292), .A2(n395), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n582), .A2(n394), .ZN(n404) );
  XNOR2_X1 U451 ( .A(n395), .B(KEYINPUT41), .ZN(n573) );
  OR2_X1 U452 ( .A1(n573), .A2(n582), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  NOR2_X1 U455 ( .A1(n398), .A2(n590), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT113), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n568), .A2(n400), .ZN(n402) );
  NAND2_X1 U458 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n405), .B(KEYINPUT48), .ZN(n539) );
  XOR2_X1 U460 ( .A(G92GAT), .B(KEYINPUT101), .Z(n407) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(n408), .B(G218GAT), .Z(n416) );
  XOR2_X1 U464 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n410) );
  XNOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT93), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n411), .B(G183GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(G169GAT), .B(G176GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n464) );
  XNOR2_X1 U470 ( .A(n464), .B(n414), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U472 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U474 ( .A(n422), .B(n421), .Z(n528) );
  INV_X1 U475 ( .A(n528), .ZN(n472) );
  NAND2_X1 U476 ( .A1(n539), .A2(n472), .ZN(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n444) );
  XOR2_X1 U479 ( .A(KEYINPUT100), .B(KEYINPUT4), .Z(n426) );
  XNOR2_X1 U480 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U482 ( .A(G57GAT), .B(KEYINPUT1), .Z(n428) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n443) );
  XOR2_X1 U486 ( .A(G113GAT), .B(KEYINPUT0), .Z(n448) );
  XOR2_X1 U487 ( .A(n431), .B(n448), .Z(n433) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U490 ( .A(G155GAT), .B(G148GAT), .Z(n435) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(G127GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U494 ( .A(G85GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U498 ( .A(n443), .B(n442), .Z(n478) );
  INV_X1 U499 ( .A(n478), .ZN(n525) );
  NAND2_X1 U500 ( .A1(n444), .A2(n525), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n581) );
  NAND2_X1 U502 ( .A1(n480), .A2(n581), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n447), .B(KEYINPUT55), .ZN(n465) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U507 ( .A(KEYINPUT65), .B(KEYINPUT91), .Z(n455) );
  NAND2_X1 U508 ( .A1(G227GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U510 ( .A(n457), .B(n456), .Z(n462) );
  XOR2_X1 U511 ( .A(KEYINPUT20), .B(KEYINPUT92), .Z(n459) );
  XNOR2_X1 U512 ( .A(G99GAT), .B(G190GAT), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT94), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U516 ( .A(n531), .ZN(n541) );
  NAND2_X1 U517 ( .A1(n465), .A2(n541), .ZN(n576) );
  NOR2_X1 U518 ( .A1(n486), .A2(n576), .ZN(n469) );
  XNOR2_X1 U519 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n467) );
  INV_X1 U520 ( .A(G190GAT), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n582), .A2(n576), .ZN(n471) );
  XNOR2_X1 U522 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n471), .B(n470), .ZN(G1348GAT) );
  NAND2_X1 U524 ( .A1(n472), .A2(n541), .ZN(n473) );
  NAND2_X1 U525 ( .A1(n480), .A2(n473), .ZN(n474) );
  XNOR2_X1 U526 ( .A(n474), .B(KEYINPUT25), .ZN(n477) );
  NOR2_X1 U527 ( .A1(n541), .A2(n480), .ZN(n475) );
  XOR2_X1 U528 ( .A(n475), .B(KEYINPUT26), .Z(n556) );
  XNOR2_X1 U529 ( .A(n528), .B(KEYINPUT27), .ZN(n481) );
  NOR2_X1 U530 ( .A1(n556), .A2(n481), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n479) );
  NOR2_X1 U532 ( .A1(n479), .A2(n478), .ZN(n485) );
  XNOR2_X1 U533 ( .A(n480), .B(KEYINPUT28), .ZN(n534) );
  INV_X1 U534 ( .A(n534), .ZN(n543) );
  XOR2_X1 U535 ( .A(KEYINPUT95), .B(n531), .Z(n482) );
  NOR2_X1 U536 ( .A1(n525), .A2(n481), .ZN(n538) );
  NAND2_X1 U537 ( .A1(n482), .A2(n538), .ZN(n483) );
  NOR2_X1 U538 ( .A1(n543), .A2(n483), .ZN(n484) );
  NOR2_X1 U539 ( .A1(n485), .A2(n484), .ZN(n500) );
  INV_X1 U540 ( .A(n486), .ZN(n552) );
  NOR2_X1 U541 ( .A1(n577), .A2(n552), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U543 ( .A1(n500), .A2(n488), .ZN(n513) );
  NOR2_X1 U544 ( .A1(n582), .A2(n395), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n489), .B(KEYINPUT78), .ZN(n503) );
  NAND2_X1 U546 ( .A1(n513), .A2(n503), .ZN(n497) );
  NOR2_X1 U547 ( .A1(n525), .A2(n497), .ZN(n490) );
  XOR2_X1 U548 ( .A(KEYINPUT34), .B(n490), .Z(n491) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n528), .A2(n497), .ZN(n492) );
  XOR2_X1 U551 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  NOR2_X1 U552 ( .A1(n497), .A2(n531), .ZN(n496) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n494) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n534), .A2(n497), .ZN(n498) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n498), .Z(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT104), .Z(n499) );
  XNOR2_X1 U560 ( .A(KEYINPUT39), .B(n499), .ZN(n506) );
  NOR2_X1 U561 ( .A1(n593), .A2(n500), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n577), .A2(n501), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT37), .B(n502), .ZN(n524) );
  NAND2_X1 U564 ( .A1(n524), .A2(n503), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT38), .B(n504), .ZN(n511) );
  NOR2_X1 U566 ( .A1(n525), .A2(n511), .ZN(n505) );
  XOR2_X1 U567 ( .A(n506), .B(n505), .Z(G1328GAT) );
  NOR2_X1 U568 ( .A1(n511), .A2(n528), .ZN(n507) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  NOR2_X1 U570 ( .A1(n511), .A2(n531), .ZN(n510) );
  XOR2_X1 U571 ( .A(G43GAT), .B(KEYINPUT106), .Z(n508) );
  XNOR2_X1 U572 ( .A(KEYINPUT40), .B(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1330GAT) );
  NOR2_X1 U574 ( .A1(n511), .A2(n534), .ZN(n512) );
  XOR2_X1 U575 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NOR2_X1 U576 ( .A1(n559), .A2(n573), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n523), .A2(n513), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n525), .A2(n520), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n520), .ZN(n517) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n531), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(n518), .Z(n519) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U587 ( .A1(n534), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n525), .A2(n533), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n533), .ZN(n532) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U600 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(KEYINPUT115), .B(n540), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n557), .A2(n541), .ZN(n542) );
  NOR2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n553), .A2(n559), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n546) );
  INV_X1 U610 ( .A(n573), .ZN(n561) );
  NAND2_X1 U611 ( .A1(n553), .A2(n561), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT116), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n550) );
  NAND2_X1 U616 ( .A1(n553), .A2(n590), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G127GAT), .B(n551), .Z(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  INV_X1 U622 ( .A(n556), .ZN(n580) );
  NAND2_X1 U623 ( .A1(n580), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT119), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n569), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n563) );
  NAND2_X1 U629 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  XOR2_X1 U632 ( .A(G155GAT), .B(KEYINPUT121), .Z(n567) );
  NAND2_X1 U633 ( .A1(n569), .A2(n590), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n572) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n573), .A2(n576), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1349GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1350GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n592) );
  NOR2_X1 U646 ( .A1(n582), .A2(n592), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n587) );
  INV_X1 U651 ( .A(n592), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n589), .A2(n395), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U654 ( .A(G204GAT), .B(n588), .Z(G1353GAT) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

