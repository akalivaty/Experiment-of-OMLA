//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(KEYINPUT2), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G113gat), .B2(G120gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G113gat), .B2(G120gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n219), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(G120gat), .ZN(new_n224));
  INV_X1    g023(.A(G113gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n223), .B(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n217), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT78), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT5), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n234), .A3(new_n216), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n226), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n216), .A4(new_n214), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n217), .B2(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n240), .A2(new_n238), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n231), .A4(new_n237), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT0), .ZN(new_n247));
  XNOR2_X1  g046(.A(G57gat), .B(G85gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n242), .A2(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT6), .B1(new_n252), .B2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT72), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(new_n261), .A3(new_n257), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT23), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(G183gat), .A3(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n282), .B(KEYINPUT64), .C1(G183gat), .C2(G190gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT66), .B(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n282), .B1(new_n291), .B2(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n274), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT28), .ZN(new_n299));
  INV_X1    g098(.A(new_n269), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n300), .A2(new_n301), .A3(new_n271), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n300), .A2(new_n301), .B1(new_n277), .B2(new_n278), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G226gat), .ZN(new_n307));
  INV_X1    g106(.A(G233gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n294), .B1(new_n287), .B2(new_n288), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI211_X1 g113(.A(KEYINPUT67), .B(new_n294), .C1(new_n287), .C2(new_n288), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n305), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n309), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n268), .B(new_n311), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n306), .A2(new_n317), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n316), .B2(new_n310), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n320), .B2(new_n268), .ZN(new_n321));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n245), .A2(KEYINPUT6), .A3(new_n250), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n254), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT37), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n320), .B2(new_n268), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n316), .A2(new_n317), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(new_n310), .B2(new_n306), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n268), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n324), .B(KEYINPUT73), .Z(new_n333));
  AOI211_X1 g132(.A(KEYINPUT38), .B(new_n333), .C1(new_n321), .C2(new_n328), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n327), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n324), .B1(new_n321), .B2(new_n328), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n328), .B2(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT38), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT31), .B(G50gat), .ZN(new_n339));
  INV_X1    g138(.A(G106gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n343));
  INV_X1    g142(.A(G228gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n308), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n234), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(new_n217), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n235), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n267), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n348), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n352), .A2(new_n356), .B1(new_n217), .B2(new_n347), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n345), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(G22gat), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT81), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n346), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n343), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G78gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n343), .B(G78gat), .C1(new_n360), .C2(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n342), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n355), .A2(G22gat), .A3(new_n359), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n364), .B2(new_n366), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT79), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G78gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n370), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n341), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n335), .A2(new_n338), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n321), .A2(KEYINPUT30), .A3(new_n324), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT75), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n321), .A2(new_n384), .A3(KEYINPUT30), .A4(new_n324), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT74), .B1(new_n321), .B2(new_n333), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n316), .A2(new_n310), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n267), .B1(new_n388), .B2(new_n319), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  INV_X1    g189(.A(new_n333), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n318), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n387), .A2(new_n392), .B1(new_n325), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n241), .A2(new_n396), .A3(new_n230), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n241), .A2(new_n230), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n228), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT39), .B1(new_n400), .B2(new_n230), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n249), .B(new_n397), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT40), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT82), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n397), .A2(new_n249), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n398), .B(KEYINPUT39), .C1(new_n230), .C2(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .A4(KEYINPUT40), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n250), .A2(new_n245), .B1(new_n402), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n381), .B1(new_n395), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g212(.A(KEYINPUT83), .B(new_n411), .C1(new_n386), .C2(new_n394), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n380), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n380), .B(new_n417), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n254), .A2(new_n326), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n395), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n373), .A2(new_n379), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT36), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n316), .A2(new_n227), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n236), .B(new_n305), .C1(new_n314), .C2(new_n315), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(G227gat), .A3(G233gat), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT70), .ZN(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n427), .A2(new_n435), .A3(new_n436), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n427), .B(KEYINPUT32), .C1(new_n436), .C2(new_n432), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n425), .A2(new_n426), .B1(G227gat), .B2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n440), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n427), .A2(new_n435), .A3(new_n436), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n428), .B(new_n433), .C1(new_n448), .C2(new_n437), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(new_n441), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n443), .B2(new_n444), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n447), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n446), .B1(new_n440), .B2(new_n442), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n441), .A3(new_n445), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n424), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n453), .B1(new_n447), .B2(new_n450), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n456), .A3(new_n452), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n423), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n454), .A2(new_n457), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n422), .A4(new_n421), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n459), .A2(new_n422), .A3(new_n460), .A4(new_n421), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n419), .A2(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n469));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(new_n472), .C1(G29gat), .C2(G36gat), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  INV_X1    g273(.A(G36gat), .ZN(new_n475));
  OAI221_X1 g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .C1(new_n470), .C2(KEYINPUT15), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n471), .B1(G29gat), .B2(G36gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT14), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT15), .B(new_n470), .C1(new_n476), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n470), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n479), .A4(new_n473), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n486), .A3(KEYINPUT87), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT87), .B1(new_n481), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n469), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(G1gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  AOI21_X1  g292(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n494), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n486), .A3(KEYINPUT17), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n489), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n487), .ZN(new_n503));
  INV_X1    g302(.A(new_n498), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n490), .A2(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n504), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n498), .A2(new_n502), .A3(new_n487), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n506), .B(KEYINPUT13), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n505), .A2(KEYINPUT18), .A3(new_n506), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G169gat), .B(G197gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT12), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(new_n514), .A3(new_n515), .A4(new_n522), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n468), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G57gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G64gat), .ZN(new_n532));
  INV_X1    g331(.A(G64gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G57gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G71gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n370), .ZN(new_n537));
  NAND2_X1  g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n535), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G71gat), .A3(G78gat), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n543), .A2(new_n545), .A3(new_n537), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n535), .A2(new_n541), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT91), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n532), .A2(new_n534), .B1(new_n540), .B2(new_n538), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n545), .A3(new_n537), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n542), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G127gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n559), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n498), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n558), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n209), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n565), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT95), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(G99gat), .A3(G106gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT8), .ZN(new_n577));
  NOR2_X1   g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n582), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  AOI21_X1  g386(.A(new_n572), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT8), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n573), .B2(KEYINPUT95), .ZN(new_n590));
  AOI211_X1 g389(.A(KEYINPUT96), .B(new_n578), .C1(new_n590), .C2(new_n576), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n582), .B1(new_n577), .B2(new_n579), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n572), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n503), .A2(new_n595), .B1(KEYINPUT41), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n490), .A2(new_n499), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(KEYINPUT93), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(KEYINPUT97), .A3(new_n605), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n571), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n570), .B2(new_n616), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n572), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n553), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(new_n588), .B2(new_n594), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n622), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n553), .A3(new_n593), .A4(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT101), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n625), .A2(new_n637), .A3(new_n628), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n625), .A2(new_n628), .A3(KEYINPUT100), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND4_X1   g441(.A1(KEYINPUT10), .A2(new_n595), .A3(new_n560), .A4(new_n561), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n631), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(KEYINPUT102), .A3(new_n631), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n632), .B(new_n635), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n631), .B(KEYINPUT103), .Z(new_n651));
  OR2_X1    g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n632), .ZN(new_n653));
  INV_X1    g452(.A(new_n635), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n621), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n530), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n420), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  INV_X1    g462(.A(new_n395), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n667), .B2(new_n665), .ZN(new_n670));
  MUX2_X1   g469(.A(new_n669), .B(new_n670), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g470(.A(new_n463), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n660), .A2(G15gat), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n458), .A2(new_n461), .ZN(new_n674));
  OAI21_X1  g473(.A(G15gat), .B1(new_n660), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(G1326gat));
  NOR3_X1   g475(.A1(new_n468), .A2(new_n529), .A3(new_n422), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n659), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n419), .A2(new_n462), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n465), .A2(new_n467), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n616), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n468), .B2(new_n617), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n656), .B(KEYINPUT105), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n526), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n571), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n687), .A2(new_n420), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G29gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n571), .A2(new_n617), .A3(new_n656), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n530), .A2(new_n474), .A3(new_n420), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(G1328gat));
  NAND4_X1  g500(.A1(new_n530), .A2(new_n475), .A3(new_n395), .A4(new_n694), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n687), .A2(new_n395), .A3(new_n691), .ZN(new_n706));
  OAI221_X1 g505(.A(new_n705), .B1(new_n703), .B2(new_n702), .C1(new_n706), .C2(new_n475), .ZN(G1329gat));
  INV_X1    g506(.A(new_n674), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n708), .A3(G43gat), .A4(new_n691), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n530), .A2(new_n463), .A3(new_n694), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(KEYINPUT47), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n712), .A2(KEYINPUT47), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(new_n422), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n684), .A2(new_n686), .A3(new_n717), .A4(new_n691), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  INV_X1    g518(.A(G50gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n677), .A2(new_n720), .A3(new_n694), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT48), .Z(G1331gat));
  AND3_X1   g522(.A1(new_n621), .A2(new_n690), .A3(new_n689), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n683), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n420), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n531), .ZN(G1332gat));
  NOR2_X1   g527(.A1(new_n725), .A2(new_n664), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  NOR3_X1   g532(.A1(new_n725), .A2(new_n672), .A3(G71gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n725), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n708), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(G71gat), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g537(.A1(new_n725), .A2(new_n422), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n370), .ZN(G1335gat));
  NAND3_X1  g539(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n616), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n468), .B2(new_n617), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n571), .A2(new_n526), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT51), .A4(new_n744), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n657), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(G85gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n420), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n571), .A2(new_n657), .A3(new_n526), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n687), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n420), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n754), .B2(new_n750), .ZN(G1336gat));
  NOR2_X1   g554(.A1(new_n664), .A2(G92gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n688), .B(new_n757), .C1(new_n747), .C2(new_n748), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n687), .A2(new_n395), .A3(new_n752), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n762));
  INV_X1    g561(.A(new_n748), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n689), .B(new_n756), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(G92gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n767), .ZN(G1337gat));
  INV_X1    g567(.A(G99gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n769), .A3(new_n463), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n753), .A2(new_n708), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n769), .ZN(G1338gat));
  NOR2_X1   g571(.A1(new_n422), .A2(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n688), .B(new_n774), .C1(new_n747), .C2(new_n748), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n687), .A2(new_n717), .A3(new_n752), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n689), .B(new_n773), .C1(new_n762), .C2(new_n763), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(G106gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(G1339gat));
  NAND3_X1  g582(.A1(new_n621), .A2(new_n690), .A3(new_n657), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n642), .A2(new_n644), .A3(new_n651), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT54), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT102), .B1(new_n648), .B2(new_n631), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n645), .A2(new_n636), .A3(new_n646), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n654), .B1(new_n652), .B2(KEYINPUT54), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n648), .B2(new_n651), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n647), .B2(new_n649), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n648), .A2(new_n651), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n635), .B1(new_n796), .B2(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n792), .A2(new_n798), .A3(new_n526), .A4(new_n650), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n505), .A2(KEYINPUT110), .A3(new_n506), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT110), .B1(new_n505), .B2(new_n506), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n800), .B(new_n801), .C1(new_n512), .C2(new_n513), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n521), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n656), .A2(new_n525), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n616), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n792), .A2(new_n650), .A3(new_n798), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n616), .A2(new_n525), .A3(new_n803), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n570), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT111), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n784), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(new_n420), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n672), .A2(new_n717), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n813), .A2(new_n664), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n225), .A3(new_n526), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n812), .A2(new_n422), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n395), .A2(new_n726), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n672), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n528), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n822), .A2(KEYINPUT112), .A3(G113gat), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT112), .B1(new_n822), .B2(G113gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n816), .B1(new_n823), .B2(new_n824), .ZN(G1340gat));
  NAND2_X1  g624(.A1(new_n656), .A2(new_n224), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT114), .Z(new_n827));
  NAND2_X1  g626(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n689), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n829), .A2(KEYINPUT113), .A3(G120gat), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n829), .B2(G120gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(G1341gat));
  INV_X1    g631(.A(new_n821), .ZN(new_n833));
  OAI21_X1  g632(.A(G127gat), .B1(new_n833), .B2(new_n570), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n815), .A2(new_n557), .A3(new_n571), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n395), .A2(new_n617), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT115), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n813), .A2(new_n837), .A3(new_n814), .A4(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(KEYINPUT117), .B2(new_n841), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(new_n845), .A3(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n817), .A2(new_n616), .A3(new_n820), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G134gat), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n844), .B(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT118), .ZN(G1343gat));
  INV_X1    g651(.A(new_n203), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n708), .A2(new_n819), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n528), .A2(new_n650), .A3(new_n798), .A4(new_n792), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n616), .B1(new_n855), .B2(new_n804), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n570), .B1(new_n856), .B2(new_n808), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n784), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n717), .A2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n812), .B2(new_n717), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(KEYINPUT119), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(KEYINPUT57), .C1(new_n812), .C2(new_n717), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n854), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n853), .B1(new_n865), .B2(new_n529), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n867));
  NAND3_X1  g666(.A1(new_n813), .A2(new_n717), .A3(new_n674), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n664), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n528), .A2(new_n205), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n866), .B(new_n867), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n526), .B(new_n854), .C1(new_n862), .C2(new_n864), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n853), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT120), .B1(new_n874), .B2(new_n853), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n868), .A2(new_n395), .A3(new_n872), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(G1344gat));
  OAI21_X1  g679(.A(new_n857), .B1(new_n658), .B2(new_n528), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n717), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n812), .A2(new_n859), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(new_n656), .A3(new_n854), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(KEYINPUT59), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n865), .B2(new_n657), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n656), .A2(new_n886), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n871), .B2(new_n891), .ZN(G1345gat));
  OAI21_X1  g691(.A(G155gat), .B1(new_n865), .B2(new_n570), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n571), .A2(new_n209), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n871), .B2(new_n894), .ZN(G1346gat));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n210), .A3(new_n839), .ZN(new_n896));
  OAI21_X1  g695(.A(G162gat), .B1(new_n865), .B2(new_n617), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NAND2_X1  g697(.A1(new_n814), .A2(new_n395), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT123), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n812), .A2(new_n726), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT124), .Z(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n526), .ZN(new_n904));
  INV_X1    g703(.A(G169gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n664), .A2(new_n420), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n463), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n817), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n529), .A2(new_n905), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n904), .A2(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  INV_X1    g709(.A(G176gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n911), .A3(new_n656), .ZN(new_n912));
  INV_X1    g711(.A(new_n908), .ZN(new_n913));
  OAI21_X1  g712(.A(G176gat), .B1(new_n913), .B2(new_n688), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(new_n297), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n902), .A2(new_n916), .A3(new_n570), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n277), .B1(new_n908), .B2(new_n571), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n919), .B(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n290), .A3(new_n616), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT61), .B(new_n278), .C1(new_n908), .C2(new_n616), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n616), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(G190gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n924), .B2(new_n927), .ZN(G1351gat));
  NAND2_X1  g727(.A1(new_n674), .A2(new_n906), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT126), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n884), .A2(G197gat), .A3(new_n528), .A4(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n708), .A2(new_n664), .A3(new_n422), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n901), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n526), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n932), .A2(new_n936), .ZN(G1352gat));
  NOR3_X1   g736(.A1(new_n934), .A2(G204gat), .A3(new_n657), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n884), .A2(new_n689), .A3(new_n930), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G204gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n259), .A3(new_n571), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n929), .A2(new_n570), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n882), .B2(new_n883), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n948), .B(new_n949), .ZN(G1354gat));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n260), .A3(new_n616), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n884), .A2(new_n616), .A3(new_n930), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n260), .ZN(G1355gat));
endmodule


