//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(new_n205), .C1(new_n206), .C2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n202), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  INV_X1    g016(.A(G127gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G134gat), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G127gat), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n217), .A2(KEYINPUT1), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G113gat), .ZN(new_n224));
  INV_X1    g023(.A(G113gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G120gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n207), .A2(new_n222), .A3(new_n215), .A4(new_n230), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n239), .A3(new_n215), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n231), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(KEYINPUT78), .A3(new_n240), .A4(new_n231), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n222), .A2(new_n230), .A3(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n216), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n233), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n252), .B(new_n235), .C1(KEYINPUT4), .C2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(KEYINPUT5), .B(new_n237), .C1(new_n246), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT79), .B1(new_n233), .B2(KEYINPUT4), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  INV_X1    g057(.A(new_n249), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT70), .B1(new_n222), .B2(new_n230), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n258), .B(new_n251), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n233), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT80), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n257), .A2(new_n261), .A3(new_n265), .A4(new_n262), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n236), .A2(KEYINPUT5), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n264), .A2(new_n245), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n255), .A2(new_n268), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n269), .A2(KEYINPUT6), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT23), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n288), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n286), .B(new_n289), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G183gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT24), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n303), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT69), .B1(new_n297), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n289), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n303), .A2(new_n307), .A3(new_n309), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n290), .A3(new_n294), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT65), .B1(new_n288), .B2(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n313), .A2(new_n314), .A3(new_n315), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n298), .ZN(new_n320));
  NAND2_X1  g119(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(G190gat), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n288), .A2(KEYINPUT23), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n302), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n322), .A2(new_n286), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n295), .A2(new_n296), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n287), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n319), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n288), .B(KEYINPUT26), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n329), .A2(new_n286), .B1(G183gat), .B2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n298), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n299), .A2(new_n301), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n331), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT28), .B1(new_n334), .B2(new_n302), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT27), .B(G183gat), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n330), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n250), .ZN(new_n342));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n343), .B(KEYINPUT64), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n250), .A2(new_n341), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n248), .A2(KEYINPUT71), .A3(new_n249), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n328), .A4(new_n339), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G71gat), .B(G99gat), .Z(new_n349));
  XNOR2_X1  g148(.A(G15gat), .B(G43gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n348), .A2(new_n357), .A3(KEYINPUT32), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n352), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n344), .B1(new_n342), .B2(new_n347), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI211_X1 g165(.A(KEYINPUT34), .B(new_n344), .C1(new_n342), .C2(new_n347), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT74), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n359), .A2(new_n368), .A3(KEYINPUT74), .A4(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  OR2_X1    g175(.A1(G197gat), .A2(G204gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT22), .ZN(new_n379));
  NAND2_X1  g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(G211gat), .A2(G218gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n380), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT76), .B1(new_n386), .B2(new_n382), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n387), .B2(new_n385), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n251), .B1(new_n391), .B2(new_n239), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n240), .A2(new_n376), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n375), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n387), .ZN(new_n397));
  INV_X1    g196(.A(new_n381), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n216), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n394), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(G22gat), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT81), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n396), .A2(new_n403), .A3(G228gat), .A4(G233gat), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n406), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n374), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n405), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n373), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n340), .A2(KEYINPUT77), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n328), .A2(new_n339), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(KEYINPUT29), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n328), .A2(new_n339), .A3(new_n429), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n393), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n328), .A2(new_n339), .A3(new_n426), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n328), .B2(new_n339), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n340), .A2(new_n430), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n393), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n424), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  INV_X1    g240(.A(new_n393), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n433), .A3(new_n423), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n444), .A3(KEYINPUT30), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n443), .A2(new_n446), .A3(new_n433), .A4(new_n423), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n445), .A2(new_n447), .B1(new_n278), .B2(new_n279), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n372), .A2(new_n420), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n412), .A2(new_n450), .A3(new_n418), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n366), .A2(new_n367), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n359), .A2(new_n452), .A3(new_n362), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n359), .B2(new_n362), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n449), .A2(KEYINPUT35), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n420), .A2(new_n448), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n266), .A2(new_n245), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n233), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n256), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n265), .B1(new_n462), .B2(new_n261), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n459), .B(new_n236), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n273), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT39), .B1(new_n234), .B2(new_n236), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n264), .A2(new_n245), .A3(new_n266), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n236), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT82), .B(new_n458), .C1(new_n465), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n236), .B1(new_n460), .B2(new_n463), .ZN(new_n471));
  INV_X1    g270(.A(new_n466), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n273), .A3(new_n464), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT82), .B1(new_n474), .B2(new_n458), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n473), .A2(KEYINPUT40), .A3(new_n273), .A4(new_n464), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n275), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n445), .A2(new_n447), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n419), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n340), .A2(new_n430), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n425), .A2(new_n427), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n429), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n482), .B(new_n433), .C1(new_n485), .C2(new_n393), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n443), .A2(new_n488), .A3(new_n482), .A4(new_n433), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n431), .A2(new_n432), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n482), .B1(new_n491), .B2(new_n442), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n441), .A2(new_n393), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n424), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n278), .A2(new_n279), .A3(new_n444), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n482), .B1(new_n443), .B2(new_n433), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n423), .B(new_n497), .C1(new_n487), .C2(new_n489), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT38), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n495), .B(new_n496), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n457), .B1(new_n481), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n453), .B2(new_n454), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT75), .B(new_n502), .C1(new_n453), .C2(new_n454), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n456), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G197gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT11), .B(G169gat), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT12), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  AOI21_X1  g318(.A(G1gat), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n518), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n525));
  AOI21_X1  g324(.A(G36gat), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n528), .B(new_n530), .C1(KEYINPUT84), .C2(new_n532), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n526), .A2(new_n527), .B1(KEYINPUT15), .B2(new_n529), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n534), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n533), .A2(new_n537), .A3(KEYINPUT17), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT17), .B1(new_n533), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n521), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n520), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n518), .A2(new_n520), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT18), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n521), .A2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n546), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n541), .B(KEYINPUT13), .Z(new_n551));
  AOI22_X1  g350(.A1(new_n547), .A2(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n546), .A4(new_n541), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n514), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n514), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n552), .A2(KEYINPUT86), .A3(new_n514), .A4(new_n553), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT87), .B1(new_n509), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n455), .A2(new_n448), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n457), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n495), .A2(new_n496), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n423), .B1(new_n487), .B2(new_n489), .ZN(new_n568));
  INV_X1    g367(.A(new_n497), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n499), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT82), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n465), .A2(new_n468), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(KEYINPUT40), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n275), .A3(new_n469), .A4(new_n476), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n420), .B1(new_n575), .B2(new_n479), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n566), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n565), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  INV_X1    g379(.A(new_n561), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n585), .A2(KEYINPUT90), .ZN(new_n586));
  NAND2_X1  g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  OR2_X1    g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(KEYINPUT90), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n587), .C1(new_n585), .C2(new_n589), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n585), .A2(KEYINPUT88), .A3(G71gat), .A4(G78gat), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n588), .B(KEYINPUT89), .Z(new_n597));
  OAI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n521), .B1(new_n584), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT91), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n203), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n600), .B(new_n602), .Z(new_n603));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n218), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n218), .B1(new_n608), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  INV_X1    g413(.A(new_n604), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n603), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n616), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n600), .B(new_n602), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT94), .B1(KEYINPUT93), .B2(KEYINPUT7), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n623), .B2(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(G85gat), .A3(G92gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G99gat), .B(G106gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n625), .A2(new_n626), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n625), .A2(new_n626), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n636), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n637), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n539), .B2(new_n538), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT97), .B1(new_n634), .B2(new_n636), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n643), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n543), .A3(new_n637), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n647), .A2(new_n649), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT98), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT92), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n220), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n204), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n538), .A2(new_n539), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n650), .A2(new_n643), .B1(new_n636), .B2(new_n634), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n652), .B(new_n653), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n648), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n655), .A2(new_n659), .B1(new_n663), .B2(new_n654), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n665), .A2(new_n663), .A3(new_n654), .A4(new_n659), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n621), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n640), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n672), .A3(new_n636), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n651), .A2(new_n605), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n661), .B2(new_n605), .ZN(new_n675));
  INV_X1    g474(.A(G230gat), .ZN(new_n676));
  INV_X1    g475(.A(G233gat), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT10), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n646), .A2(new_n680), .A3(new_n598), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n675), .B2(KEYINPUT10), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n598), .B1(new_n650), .B2(new_n643), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n646), .A2(new_n598), .B1(new_n684), .B2(new_n673), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(KEYINPUT100), .A3(new_n680), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n681), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n679), .B1(new_n687), .B2(new_n678), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n681), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n685), .B2(new_n680), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n646), .A2(new_n598), .ZN(new_n696));
  AND4_X1   g495(.A1(KEYINPUT100), .A2(new_n696), .A3(new_n680), .A4(new_n674), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n678), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n679), .A3(new_n691), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n693), .A2(new_n701), .A3(KEYINPUT101), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n669), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT102), .B1(new_n583), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n706), .C1(new_n562), .C2(new_n582), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n281), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g511(.A(KEYINPUT16), .B(G8gat), .Z(new_n713));
  OAI211_X1 g512(.A(new_n480), .B(new_n713), .C1(new_n708), .C2(new_n710), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n509), .A2(KEYINPUT87), .A3(new_n561), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n580), .B1(new_n579), .B2(new_n581), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n707), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n709), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n583), .A2(KEYINPUT102), .A3(new_n707), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n479), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n714), .B1(new_n720), .B2(new_n517), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1325gat));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n453), .A2(new_n454), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(G15gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n708), .B2(new_n710), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n508), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n505), .A2(new_n507), .A3(KEYINPUT103), .A4(new_n506), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n718), .B2(new_n719), .ZN(new_n735));
  INV_X1    g534(.A(G15gat), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n726), .B(new_n730), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n734), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n708), .B2(new_n710), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G15gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n726), .B1(new_n741), .B2(new_n730), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n738), .A2(new_n742), .ZN(G1326gat));
  OAI21_X1  g542(.A(new_n419), .B1(new_n708), .B2(new_n710), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT43), .B(G22gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1327gat));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n704), .A2(new_n705), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n668), .A3(new_n621), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n562), .B2(new_n582), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n281), .A2(new_n523), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n667), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n579), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n621), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n748), .A2(new_n561), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n732), .A2(new_n501), .A3(new_n733), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n667), .B1(new_n760), .B2(new_n565), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n757), .B(new_n759), .C1(new_n761), .C2(KEYINPUT44), .ZN(new_n762));
  OAI21_X1  g561(.A(G29gat), .B1(new_n762), .B2(new_n280), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n751), .A2(KEYINPUT45), .A3(new_n523), .A4(new_n281), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n754), .A2(new_n763), .A3(new_n764), .ZN(G1328gat));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n479), .A2(G36gat), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n751), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n751), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n762), .B2(new_n479), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G36gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n762), .A2(new_n771), .A3(new_n479), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT106), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n770), .B(new_n777), .C1(new_n773), .C2(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1329gat));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n565), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n668), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n781), .A2(new_n755), .B1(new_n579), .B2(new_n756), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(G43gat), .A3(new_n739), .A4(new_n759), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n752), .A2(new_n728), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n783), .B(new_n785), .C1(new_n786), .C2(G43gat), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1330gat));
  OAI21_X1  g588(.A(G50gat), .B1(new_n762), .B2(new_n420), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n420), .A2(G50gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n752), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT48), .Z(G1331gat));
  AND4_X1   g592(.A1(new_n561), .A2(new_n780), .A3(new_n669), .A4(new_n748), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n281), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g595(.A(new_n479), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT108), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1333gat));
  XNOR2_X1  g600(.A(new_n727), .B(KEYINPUT109), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(G71gat), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n739), .A2(G71gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1334gat));
  NAND2_X1  g607(.A1(new_n794), .A2(new_n419), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n761), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n758), .A2(new_n581), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n761), .A2(new_n811), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n813), .A4(new_n812), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n280), .A2(G85gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n816), .A2(new_n748), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n813), .A2(new_n748), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n782), .A2(new_n822), .A3(new_n281), .A4(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n757), .B(new_n823), .C1(new_n761), .C2(KEYINPUT44), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT110), .B1(new_n825), .B2(new_n280), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(G85gat), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n821), .A2(new_n827), .A3(KEYINPUT112), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1336gat));
  INV_X1    g631(.A(new_n825), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n624), .B1(new_n833), .B2(new_n480), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n479), .A2(G92gat), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n816), .A2(new_n748), .A3(new_n819), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n814), .B2(new_n815), .ZN(new_n840));
  INV_X1    g639(.A(new_n839), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n817), .A2(new_n813), .A3(new_n812), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n749), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n834), .B1(new_n843), .B2(new_n836), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(G1337gat));
  NAND3_X1  g645(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n739), .ZN(new_n847));
  XNOR2_X1  g646(.A(KEYINPUT115), .B(G99gat), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n825), .B2(new_n734), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n728), .A2(new_n848), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n816), .A2(new_n748), .A3(new_n819), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1338gat));
  INV_X1    g653(.A(G106gat), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n833), .B2(new_n419), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n420), .A2(G106gat), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n816), .A2(new_n748), .A3(new_n819), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n843), .B2(new_n858), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(G1339gat));
  NOR2_X1   g662(.A1(new_n687), .A2(new_n678), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n691), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n687), .A2(new_n678), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n700), .A2(new_n867), .A3(KEYINPUT54), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT55), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n550), .A2(new_n551), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n540), .A2(new_n546), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(G229gat), .A3(G233gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n559), .A2(new_n560), .B1(new_n513), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n701), .B1(new_n874), .B2(new_n667), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n667), .A2(new_n561), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n869), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n698), .A2(new_n865), .A3(new_n699), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n687), .B2(new_n678), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n699), .B(new_n681), .C1(new_n683), .C2(new_n686), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n692), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT55), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n866), .A2(new_n868), .A3(KEYINPUT116), .A4(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n874), .A2(new_n667), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n877), .A2(new_n886), .B1(new_n748), .B2(new_n887), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n888), .A2(new_n758), .B1(new_n581), .B2(new_n706), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n480), .A2(new_n280), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n727), .A2(new_n889), .A3(new_n420), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n225), .B1(new_n891), .B2(new_n581), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT117), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n372), .A2(new_n420), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n889), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n225), .A3(new_n581), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n897), .ZN(G1340gat));
  AOI21_X1  g697(.A(G120gat), .B1(new_n896), .B2(new_n748), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n749), .A2(new_n223), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n891), .B2(new_n900), .ZN(G1341gat));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n218), .A3(new_n758), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n891), .A2(new_n758), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n218), .ZN(G1342gat));
  NAND2_X1  g703(.A1(new_n891), .A2(new_n668), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G134gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n896), .A2(new_n220), .A3(new_n668), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n910));
  OAI221_X1 g709(.A(new_n906), .B1(KEYINPUT56), .B2(new_n907), .C1(new_n909), .C2(new_n910), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n734), .A2(new_n890), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n561), .A2(G141gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n913), .A2(new_n419), .A3(new_n889), .A4(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(KEYINPUT120), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n877), .A2(new_n886), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n748), .A2(new_n887), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n758), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n706), .A2(new_n581), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n918), .B1(new_n923), .B2(new_n420), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n419), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n912), .B(KEYINPUT119), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n581), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n917), .B1(new_n928), .B2(G141gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(KEYINPUT58), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n929), .B(new_n931), .ZN(G1344gat));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(KEYINPUT121), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n926), .A2(new_n927), .ZN(new_n935));
  OAI211_X1 g734(.A(G148gat), .B(new_n934), .C1(new_n935), .C2(new_n749), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n923), .A2(new_n912), .A3(new_n420), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n210), .A3(new_n748), .ZN(new_n938));
  INV_X1    g737(.A(new_n935), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n210), .B1(new_n939), .B2(new_n748), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n941));
  OAI211_X1 g740(.A(new_n936), .B(new_n938), .C1(new_n940), .C2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n935), .B2(new_n621), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n203), .A3(new_n758), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  AOI21_X1  g744(.A(G162gat), .B1(new_n937), .B2(new_n668), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n667), .A2(new_n204), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n939), .B2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n281), .A2(new_n479), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n889), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n895), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n291), .A3(new_n581), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n802), .A2(new_n419), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n949), .B(new_n954), .C1(new_n921), .C2(new_n922), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n889), .A2(KEYINPUT122), .A3(new_n949), .A4(new_n954), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n581), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(G169gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n959), .B2(G169gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n953), .B1(new_n961), .B2(new_n962), .ZN(G1348gat));
  NOR2_X1   g762(.A1(new_n749), .A2(new_n292), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n957), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n292), .B1(new_n951), .B2(new_n749), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n957), .A2(KEYINPUT124), .A3(new_n958), .A4(new_n964), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT125), .ZN(G1349gat));
  NAND3_X1  g770(.A1(new_n957), .A2(new_n758), .A3(new_n958), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n333), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n958), .A4(new_n758), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n952), .A2(new_n337), .A3(new_n758), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT60), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n981), .A3(new_n978), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n952), .A2(new_n302), .A3(new_n668), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n957), .A2(new_n668), .A3(new_n958), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(G190gat), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n985), .B2(G190gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G1351gat));
  NAND2_X1  g788(.A1(new_n734), .A2(new_n949), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n923), .A2(new_n990), .A3(new_n420), .ZN(new_n991));
  AOI21_X1  g790(.A(G197gat), .B1(new_n991), .B2(new_n581), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n990), .B1(new_n924), .B2(new_n925), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n581), .A2(G197gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G1352gat));
  INV_X1    g794(.A(new_n991), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n996), .A2(G204gat), .A3(new_n749), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n993), .A2(new_n748), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G204gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n1000), .ZN(G1353gat));
  OR3_X1    g800(.A1(new_n996), .A2(G211gat), .A3(new_n621), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n993), .A2(new_n758), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  INV_X1    g805(.A(G218gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n993), .B2(new_n668), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n996), .A2(G218gat), .A3(new_n667), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1010));
  OR3_X1    g809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


