

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725;

  INV_X1 U367 ( .A(G953), .ZN(n711) );
  XNOR2_X1 U368 ( .A(n455), .B(n454), .ZN(n569) );
  NAND2_X1 U369 ( .A1(n652), .A2(n653), .ZN(n649) );
  XNOR2_X2 U370 ( .A(n536), .B(KEYINPUT1), .ZN(n650) );
  XNOR2_X2 U371 ( .A(G122), .B(G104), .ZN(n389) );
  INV_X2 U372 ( .A(n389), .ZN(n505) );
  XNOR2_X2 U373 ( .A(n346), .B(n521), .ZN(n722) );
  AND2_X2 U374 ( .A1(n547), .A2(n394), .ZN(n346) );
  NOR2_X2 U375 ( .A1(n724), .A2(n725), .ZN(n590) );
  NOR2_X1 U376 ( .A1(n650), .A2(n649), .ZN(n540) );
  INV_X2 U377 ( .A(n569), .ZN(n652) );
  AND2_X1 U378 ( .A1(n359), .A2(n358), .ZN(n686) );
  AND2_X2 U379 ( .A1(n413), .A2(n344), .ZN(n692) );
  XNOR2_X1 U380 ( .A(n407), .B(n528), .ZN(n721) );
  NAND2_X1 U381 ( .A1(n527), .A2(n571), .ZN(n407) );
  XNOR2_X1 U382 ( .A(n580), .B(KEYINPUT38), .ZN(n639) );
  NAND2_X2 U383 ( .A1(n368), .A2(n369), .ZN(n656) );
  XNOR2_X1 U384 ( .A(n495), .B(n456), .ZN(n375) );
  XNOR2_X1 U385 ( .A(n435), .B(G128), .ZN(n495) );
  INV_X1 U386 ( .A(KEYINPUT71), .ZN(n388) );
  NOR2_X1 U387 ( .A1(n529), .A2(n556), .ZN(n547) );
  XNOR2_X1 U388 ( .A(n707), .B(G146), .ZN(n473) );
  NAND2_X2 U389 ( .A1(n373), .A2(n414), .ZN(n710) );
  NOR2_X1 U390 ( .A1(n632), .A2(n415), .ZN(n414) );
  XNOR2_X1 U391 ( .A(n364), .B(n374), .ZN(n373) );
  INV_X1 U392 ( .A(n719), .ZN(n415) );
  XNOR2_X1 U393 ( .A(n375), .B(n437), .ZN(n707) );
  XOR2_X1 U394 ( .A(G137), .B(G134), .Z(n437) );
  NAND2_X1 U395 ( .A1(n656), .A2(n640), .ZN(n566) );
  XNOR2_X1 U396 ( .A(n517), .B(n516), .ZN(n532) );
  XNOR2_X1 U397 ( .A(n515), .B(G475), .ZN(n516) );
  NOR2_X1 U398 ( .A1(G902), .A2(n682), .ZN(n517) );
  XNOR2_X1 U399 ( .A(n463), .B(n462), .ZN(n536) );
  XNOR2_X1 U400 ( .A(n656), .B(n376), .ZN(n556) );
  INV_X1 U401 ( .A(KEYINPUT6), .ZN(n376) );
  NOR2_X1 U402 ( .A1(n710), .A2(n634), .ZN(n408) );
  INV_X1 U403 ( .A(KEYINPUT0), .ZN(n362) );
  XOR2_X1 U404 ( .A(G125), .B(G146), .Z(n478) );
  NAND2_X1 U405 ( .A1(G234), .A2(G237), .ZN(n490) );
  XNOR2_X1 U406 ( .A(G116), .B(G131), .ZN(n467) );
  INV_X1 U407 ( .A(KEYINPUT91), .ZN(n466) );
  XNOR2_X1 U408 ( .A(n478), .B(n411), .ZN(n512) );
  INV_X1 U409 ( .A(KEYINPUT10), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n386), .B(n482), .ZN(n600) );
  XNOR2_X1 U411 ( .A(n392), .B(n480), .ZN(n482) );
  XNOR2_X1 U412 ( .A(n701), .B(n477), .ZN(n386) );
  INV_X1 U413 ( .A(n570), .ZN(n418) );
  XNOR2_X1 U414 ( .A(G119), .B(G110), .ZN(n446) );
  XOR2_X1 U415 ( .A(KEYINPUT74), .B(G140), .Z(n447) );
  XNOR2_X1 U416 ( .A(n512), .B(n409), .ZN(n444) );
  XNOR2_X1 U417 ( .A(n442), .B(n410), .ZN(n409) );
  INV_X1 U418 ( .A(KEYINPUT24), .ZN(n410) );
  XNOR2_X1 U419 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U420 ( .A(n473), .B(n391), .ZN(n674) );
  XNOR2_X1 U421 ( .A(n458), .B(n461), .ZN(n391) );
  XNOR2_X1 U422 ( .A(n460), .B(n459), .ZN(n461) );
  AND2_X1 U423 ( .A1(n347), .A2(n433), .ZN(n431) );
  XNOR2_X1 U424 ( .A(n582), .B(KEYINPUT70), .ZN(n583) );
  XNOR2_X1 U425 ( .A(n557), .B(KEYINPUT102), .ZN(n564) );
  XNOR2_X1 U426 ( .A(n422), .B(KEYINPUT22), .ZN(n529) );
  OR2_X1 U427 ( .A1(n604), .A2(n370), .ZN(n369) );
  AND2_X1 U428 ( .A1(n367), .A2(n348), .ZN(n368) );
  NAND2_X1 U429 ( .A1(n372), .A2(n371), .ZN(n370) );
  BUF_X1 U430 ( .A(n536), .Z(n401) );
  NAND2_X1 U431 ( .A1(n599), .A2(n598), .ZN(n413) );
  NAND2_X1 U432 ( .A1(n692), .A2(G475), .ZN(n412) );
  NOR2_X1 U433 ( .A1(n425), .A2(n429), .ZN(n424) );
  NAND2_X1 U434 ( .A1(n430), .A2(n711), .ZN(n429) );
  NOR2_X1 U435 ( .A1(n344), .A2(n426), .ZN(n425) );
  OR2_X1 U436 ( .A1(n347), .A2(n433), .ZN(n430) );
  XNOR2_X1 U437 ( .A(n637), .B(KEYINPUT79), .ZN(n638) );
  NOR2_X1 U438 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U439 ( .A1(n344), .A2(KEYINPUT116), .ZN(n423) );
  NOR2_X1 U440 ( .A1(G953), .A2(G237), .ZN(n508) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(G110), .Z(n476) );
  XNOR2_X1 U442 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n456) );
  XNOR2_X1 U443 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  XNOR2_X1 U444 ( .A(n479), .B(n481), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n478), .B(n345), .ZN(n479) );
  AND2_X1 U446 ( .A1(G953), .A2(G902), .ZN(n492) );
  XNOR2_X1 U447 ( .A(n507), .B(n356), .ZN(n509) );
  XNOR2_X1 U448 ( .A(G113), .B(KEYINPUT95), .ZN(n507) );
  XNOR2_X1 U449 ( .A(n357), .B(KEYINPUT94), .ZN(n356) );
  INV_X1 U450 ( .A(KEYINPUT11), .ZN(n357) );
  XNOR2_X1 U451 ( .A(n476), .B(n439), .ZN(n457) );
  XOR2_X1 U452 ( .A(G107), .B(G104), .Z(n439) );
  XOR2_X1 U453 ( .A(G131), .B(G140), .Z(n513) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n666) );
  INV_X1 U455 ( .A(KEYINPUT52), .ZN(n397) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n374) );
  XOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .Z(n594) );
  NOR2_X1 U458 ( .A1(G902), .A2(G237), .ZN(n483) );
  INV_X1 U459 ( .A(G902), .ZN(n371) );
  INV_X1 U460 ( .A(G472), .ZN(n372) );
  XNOR2_X1 U461 ( .A(n473), .B(n474), .ZN(n604) );
  XNOR2_X1 U462 ( .A(n385), .B(n496), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n505), .B(n387), .ZN(n385) );
  XNOR2_X1 U464 ( .A(n388), .B(KEYINPUT16), .ZN(n387) );
  XOR2_X1 U465 ( .A(G116), .B(G107), .Z(n496) );
  NOR2_X1 U466 ( .A1(n568), .A2(n416), .ZN(n581) );
  NAND2_X1 U467 ( .A1(n652), .A2(n417), .ZN(n416) );
  NOR2_X1 U468 ( .A1(n401), .A2(n418), .ZN(n417) );
  NOR2_X1 U469 ( .A1(n401), .A2(n577), .ZN(n588) );
  XNOR2_X1 U470 ( .A(G128), .B(G137), .ZN(n443) );
  XNOR2_X1 U471 ( .A(n379), .B(n353), .ZN(n378) );
  NAND2_X1 U472 ( .A1(n692), .A2(G210), .ZN(n379) );
  XNOR2_X1 U473 ( .A(n560), .B(n393), .ZN(n561) );
  XNOR2_X1 U474 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n393) );
  AND2_X1 U475 ( .A1(n380), .A2(n558), .ZN(n629) );
  XNOR2_X1 U476 ( .A(n381), .B(KEYINPUT36), .ZN(n380) );
  NOR2_X1 U477 ( .A1(n564), .A2(n563), .ZN(n381) );
  NOR2_X1 U478 ( .A1(n650), .A2(n652), .ZN(n394) );
  NAND2_X1 U479 ( .A1(n530), .A2(n569), .ZN(n615) );
  XNOR2_X1 U480 ( .A(n384), .B(n383), .ZN(n530) );
  INV_X1 U481 ( .A(KEYINPUT65), .ZN(n383) );
  NOR2_X1 U482 ( .A1(n529), .A2(n351), .ZN(n384) );
  XNOR2_X1 U483 ( .A(n360), .B(KEYINPUT98), .ZN(n627) );
  AND2_X1 U484 ( .A1(n539), .A2(n361), .ZN(n611) );
  NOR2_X1 U485 ( .A1(n401), .A2(n656), .ZN(n361) );
  XNOR2_X1 U486 ( .A(n412), .B(n685), .ZN(n359) );
  XNOR2_X1 U487 ( .A(n673), .B(n404), .ZN(n678) );
  NOR2_X1 U488 ( .A1(n638), .A2(n423), .ZN(n432) );
  NAND2_X1 U489 ( .A1(n382), .A2(n408), .ZN(n344) );
  AND2_X1 U490 ( .A1(G224), .A2(n711), .ZN(n345) );
  AND2_X1 U491 ( .A1(n671), .A2(n670), .ZN(n347) );
  NAND2_X1 U492 ( .A1(G902), .A2(G472), .ZN(n348) );
  NOR2_X1 U493 ( .A1(n546), .A2(n419), .ZN(n349) );
  INV_X1 U494 ( .A(n656), .ZN(n574) );
  OR2_X1 U495 ( .A1(n551), .A2(n494), .ZN(n350) );
  OR2_X1 U496 ( .A1(n558), .A2(n656), .ZN(n351) );
  XNOR2_X1 U497 ( .A(n488), .B(KEYINPUT19), .ZN(n489) );
  XOR2_X1 U498 ( .A(KEYINPUT85), .B(n441), .Z(n696) );
  INV_X1 U499 ( .A(n696), .ZN(n358) );
  XNOR2_X1 U500 ( .A(n605), .B(KEYINPUT62), .ZN(n352) );
  XOR2_X1 U501 ( .A(n602), .B(n601), .Z(n353) );
  XOR2_X1 U502 ( .A(KEYINPUT81), .B(KEYINPUT45), .Z(n354) );
  XOR2_X1 U503 ( .A(n603), .B(KEYINPUT56), .Z(n355) );
  INV_X1 U504 ( .A(KEYINPUT116), .ZN(n433) );
  XNOR2_X1 U505 ( .A(n541), .B(KEYINPUT88), .ZN(n537) );
  XNOR2_X2 U506 ( .A(n363), .B(n362), .ZN(n541) );
  NOR2_X1 U507 ( .A1(n533), .A2(n534), .ZN(n360) );
  NOR2_X1 U508 ( .A1(n545), .A2(n644), .ZN(n546) );
  INV_X1 U509 ( .A(n607), .ZN(n419) );
  NAND2_X2 U510 ( .A1(n578), .A2(n350), .ZN(n363) );
  NAND2_X1 U511 ( .A1(n366), .A2(n365), .ZN(n364) );
  XNOR2_X1 U512 ( .A(n590), .B(KEYINPUT46), .ZN(n365) );
  AND2_X1 U513 ( .A1(n591), .A2(n395), .ZN(n366) );
  NAND2_X1 U514 ( .A1(n604), .A2(G472), .ZN(n367) );
  XNOR2_X1 U515 ( .A(n375), .B(n434), .ZN(n480) );
  XNOR2_X1 U516 ( .A(n377), .B(n355), .ZN(G51) );
  NAND2_X1 U517 ( .A1(n378), .A2(n358), .ZN(n377) );
  NOR2_X1 U518 ( .A1(n382), .A2(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U519 ( .A1(n382), .A2(n711), .ZN(n700) );
  NAND2_X1 U520 ( .A1(n596), .A2(n382), .ZN(n599) );
  XNOR2_X2 U521 ( .A(n400), .B(n354), .ZN(n382) );
  XNOR2_X2 U522 ( .A(n562), .B(n489), .ZN(n578) );
  NAND2_X1 U523 ( .A1(n565), .A2(n640), .ZN(n562) );
  NOR2_X2 U524 ( .A1(n600), .A2(n594), .ZN(n485) );
  NAND2_X1 U525 ( .A1(n390), .A2(n406), .ZN(n531) );
  NOR2_X1 U526 ( .A1(n405), .A2(n722), .ZN(n390) );
  NAND2_X1 U527 ( .A1(n541), .A2(n520), .ZN(n422) );
  XNOR2_X1 U528 ( .A(n525), .B(n524), .ZN(n527) );
  NAND2_X1 U529 ( .A1(n427), .A2(n424), .ZN(n428) );
  NAND2_X1 U530 ( .A1(n662), .A2(n588), .ZN(n589) );
  XNOR2_X2 U531 ( .A(n587), .B(KEYINPUT41), .ZN(n662) );
  INV_X1 U532 ( .A(n629), .ZN(n395) );
  XNOR2_X1 U533 ( .A(n396), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U534 ( .A1(n402), .A2(n358), .ZN(n396) );
  NOR2_X2 U535 ( .A1(n432), .A2(n428), .ZN(n672) );
  NAND2_X1 U536 ( .A1(n665), .A2(n664), .ZN(n398) );
  NAND2_X1 U537 ( .A1(n399), .A2(n646), .ZN(n647) );
  XNOR2_X1 U538 ( .A(n645), .B(KEYINPUT113), .ZN(n399) );
  NAND2_X1 U539 ( .A1(n669), .A2(n537), .ZN(n525) );
  XNOR2_X2 U540 ( .A(n523), .B(KEYINPUT33), .ZN(n669) );
  NAND2_X1 U541 ( .A1(n420), .A2(n349), .ZN(n400) );
  XNOR2_X1 U542 ( .A(n606), .B(n352), .ZN(n402) );
  XNOR2_X2 U543 ( .A(n403), .B(n475), .ZN(n701) );
  INV_X1 U544 ( .A(G143), .ZN(n435) );
  INV_X1 U545 ( .A(n674), .ZN(n404) );
  INV_X1 U546 ( .A(n615), .ZN(n405) );
  INV_X1 U547 ( .A(n721), .ZN(n406) );
  NAND2_X1 U548 ( .A1(n581), .A2(n639), .ZN(n584) );
  XNOR2_X1 U549 ( .A(n449), .B(n450), .ZN(n691) );
  XNOR2_X2 U550 ( .A(n485), .B(n484), .ZN(n565) );
  XNOR2_X1 U551 ( .A(n531), .B(n421), .ZN(n420) );
  INV_X1 U552 ( .A(KEYINPUT44), .ZN(n421) );
  NAND2_X1 U553 ( .A1(n638), .A2(n431), .ZN(n427) );
  INV_X1 U554 ( .A(n431), .ZN(n426) );
  XOR2_X1 U555 ( .A(n447), .B(n446), .Z(n436) );
  AND2_X1 U556 ( .A1(n508), .A2(G214), .ZN(n438) );
  XOR2_X1 U557 ( .A(KEYINPUT47), .B(n579), .Z(n440) );
  XNOR2_X1 U558 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U559 ( .A(n469), .B(n468), .ZN(n472) );
  XNOR2_X1 U560 ( .A(n472), .B(n475), .ZN(n474) );
  XNOR2_X1 U561 ( .A(n509), .B(n438), .ZN(n510) );
  XNOR2_X1 U562 ( .A(n457), .B(n513), .ZN(n458) );
  INV_X1 U563 ( .A(KEYINPUT39), .ZN(n582) );
  XNOR2_X1 U564 ( .A(n448), .B(n436), .ZN(n449) );
  INV_X1 U565 ( .A(KEYINPUT34), .ZN(n524) );
  XNOR2_X1 U566 ( .A(n584), .B(n583), .ZN(n592) );
  INV_X1 U567 ( .A(KEYINPUT117), .ZN(n603) );
  NOR2_X1 U568 ( .A1(G952), .A2(n711), .ZN(n441) );
  XNOR2_X1 U569 ( .A(n444), .B(n443), .ZN(n450) );
  NAND2_X1 U570 ( .A1(G234), .A2(n711), .ZN(n445) );
  XOR2_X1 U571 ( .A(KEYINPUT8), .B(n445), .Z(n499) );
  NAND2_X1 U572 ( .A1(G221), .A2(n499), .ZN(n448) );
  NOR2_X1 U573 ( .A1(n691), .A2(G902), .ZN(n455) );
  XOR2_X1 U574 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n453) );
  INV_X1 U575 ( .A(n594), .ZN(n597) );
  NAND2_X1 U576 ( .A1(G234), .A2(n597), .ZN(n451) );
  XNOR2_X1 U577 ( .A(KEYINPUT20), .B(n451), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n518), .A2(G217), .ZN(n452) );
  XNOR2_X1 U579 ( .A(n453), .B(n452), .ZN(n454) );
  AND2_X1 U580 ( .A1(G227), .A2(n711), .ZN(n460) );
  XOR2_X1 U581 ( .A(G101), .B(KEYINPUT75), .Z(n459) );
  NOR2_X1 U582 ( .A1(G902), .A2(n674), .ZN(n463) );
  XNOR2_X1 U583 ( .A(KEYINPUT68), .B(G469), .ZN(n462) );
  INV_X1 U584 ( .A(n650), .ZN(n558) );
  XOR2_X1 U585 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n465) );
  NAND2_X1 U586 ( .A1(n508), .A2(G210), .ZN(n464) );
  XNOR2_X1 U587 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U588 ( .A(G101), .B(G119), .Z(n471) );
  XNOR2_X1 U589 ( .A(G113), .B(KEYINPUT3), .ZN(n470) );
  XNOR2_X1 U590 ( .A(n471), .B(n470), .ZN(n475) );
  XNOR2_X1 U591 ( .A(n476), .B(KEYINPUT76), .ZN(n477) );
  INV_X1 U592 ( .A(KEYINPUT83), .ZN(n481) );
  XOR2_X1 U593 ( .A(KEYINPUT72), .B(n483), .Z(n486) );
  NAND2_X1 U594 ( .A1(G210), .A2(n486), .ZN(n484) );
  NAND2_X1 U595 ( .A1(G214), .A2(n486), .ZN(n487) );
  XNOR2_X1 U596 ( .A(n487), .B(KEYINPUT86), .ZN(n640) );
  INV_X1 U597 ( .A(KEYINPUT67), .ZN(n488) );
  XNOR2_X1 U598 ( .A(KEYINPUT14), .B(n490), .ZN(n493) );
  NAND2_X1 U599 ( .A1(G952), .A2(n493), .ZN(n491) );
  XOR2_X1 U600 ( .A(KEYINPUT87), .B(n491), .Z(n667) );
  NOR2_X1 U601 ( .A1(G953), .A2(n667), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n493), .A2(n492), .ZN(n549) );
  NOR2_X1 U603 ( .A1(G898), .A2(n549), .ZN(n494) );
  XOR2_X1 U604 ( .A(n495), .B(G134), .Z(n498) );
  XNOR2_X1 U605 ( .A(n496), .B(G122), .ZN(n497) );
  XNOR2_X1 U606 ( .A(n498), .B(n497), .ZN(n503) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n501) );
  NAND2_X1 U608 ( .A1(G217), .A2(n499), .ZN(n500) );
  XNOR2_X1 U609 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n503), .B(n502), .ZN(n687) );
  NOR2_X1 U611 ( .A1(n687), .A2(G902), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n504), .B(G478), .ZN(n534) );
  INV_X1 U613 ( .A(n534), .ZN(n526) );
  XNOR2_X1 U614 ( .A(n505), .B(G143), .ZN(n506) );
  XNOR2_X1 U615 ( .A(n506), .B(KEYINPUT12), .ZN(n511) );
  XNOR2_X1 U616 ( .A(n511), .B(n510), .ZN(n514) );
  XNOR2_X1 U617 ( .A(n513), .B(n512), .ZN(n708) );
  XNOR2_X1 U618 ( .A(n514), .B(n708), .ZN(n682) );
  XNOR2_X1 U619 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n515) );
  NOR2_X1 U620 ( .A1(n526), .A2(n532), .ZN(n641) );
  NAND2_X1 U621 ( .A1(n518), .A2(G221), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n519), .B(KEYINPUT21), .ZN(n554) );
  INV_X1 U623 ( .A(n554), .ZN(n653) );
  AND2_X1 U624 ( .A1(n641), .A2(n653), .ZN(n520) );
  XNOR2_X1 U625 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n521) );
  XNOR2_X1 U626 ( .A(n540), .B(KEYINPUT100), .ZN(n522) );
  NAND2_X1 U627 ( .A1(n522), .A2(n556), .ZN(n523) );
  AND2_X1 U628 ( .A1(n532), .A2(n526), .ZN(n571) );
  XOR2_X1 U629 ( .A(KEYINPUT35), .B(KEYINPUT77), .Z(n528) );
  XOR2_X1 U630 ( .A(n532), .B(KEYINPUT97), .Z(n533) );
  NAND2_X1 U631 ( .A1(n534), .A2(n533), .ZN(n622) );
  INV_X1 U632 ( .A(n627), .ZN(n617) );
  NAND2_X1 U633 ( .A1(n622), .A2(n617), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(KEYINPUT99), .ZN(n644) );
  INV_X1 U635 ( .A(n537), .ZN(n538) );
  NOR2_X1 U636 ( .A1(n649), .A2(n538), .ZN(n539) );
  XOR2_X1 U637 ( .A(KEYINPUT31), .B(KEYINPUT93), .Z(n544) );
  NAND2_X1 U638 ( .A1(n656), .A2(n540), .ZN(n659) );
  INV_X1 U639 ( .A(n659), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U641 ( .A(n544), .B(n543), .ZN(n626) );
  NOR2_X1 U642 ( .A1(n611), .A2(n626), .ZN(n545) );
  AND2_X1 U643 ( .A1(n650), .A2(n547), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n652), .A2(n548), .ZN(n607) );
  XOR2_X1 U645 ( .A(n549), .B(KEYINPUT101), .Z(n550) );
  NOR2_X1 U646 ( .A1(G900), .A2(n550), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U648 ( .A1(n554), .A2(n553), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n573) );
  NOR2_X1 U650 ( .A1(n622), .A2(n573), .ZN(n555) );
  NAND2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U652 ( .A1(n558), .A2(n564), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n640), .A2(n559), .ZN(n560) );
  NOR2_X1 U654 ( .A1(n565), .A2(n561), .ZN(n632) );
  BUF_X1 U655 ( .A(n562), .Z(n563) );
  INV_X1 U656 ( .A(n565), .ZN(n580) );
  XOR2_X1 U657 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n567) );
  XOR2_X1 U658 ( .A(n567), .B(n566), .Z(n568) );
  NAND2_X1 U659 ( .A1(n581), .A2(n571), .ZN(n572) );
  NOR2_X1 U660 ( .A1(n580), .A2(n572), .ZN(n620) );
  NOR2_X1 U661 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U662 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n575) );
  XNOR2_X1 U663 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n588), .A2(n578), .ZN(n621) );
  NOR2_X1 U665 ( .A1(n621), .A2(n644), .ZN(n579) );
  NOR2_X1 U666 ( .A1(n620), .A2(n440), .ZN(n591) );
  NOR2_X1 U667 ( .A1(n592), .A2(n622), .ZN(n585) );
  XNOR2_X1 U668 ( .A(n585), .B(KEYINPUT40), .ZN(n724) );
  NAND2_X1 U669 ( .A1(n639), .A2(n640), .ZN(n643) );
  INV_X1 U670 ( .A(n643), .ZN(n586) );
  NAND2_X1 U671 ( .A1(n586), .A2(n641), .ZN(n587) );
  XOR2_X1 U672 ( .A(KEYINPUT42), .B(n589), .Z(n725) );
  OR2_X1 U673 ( .A1(n592), .A2(n617), .ZN(n593) );
  XNOR2_X1 U674 ( .A(KEYINPUT106), .B(n593), .ZN(n719) );
  XNOR2_X1 U675 ( .A(n710), .B(KEYINPUT73), .ZN(n595) );
  AND2_X1 U676 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n634) );
  OR2_X1 U678 ( .A1(n597), .A2(n634), .ZN(n598) );
  XOR2_X1 U679 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n602) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT82), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n692), .A2(G472), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT107), .ZN(n605) );
  XNOR2_X1 U683 ( .A(G101), .B(KEYINPUT108), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(n607), .ZN(G3) );
  XOR2_X1 U685 ( .A(G104), .B(KEYINPUT109), .Z(n610) );
  INV_X1 U686 ( .A(n622), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n611), .A2(n624), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n610), .B(n609), .ZN(G6) );
  XOR2_X1 U689 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U690 ( .A1(n611), .A2(n627), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U692 ( .A(G107), .B(n614), .ZN(G9) );
  XNOR2_X1 U693 ( .A(G110), .B(KEYINPUT110), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n616), .B(n615), .ZN(G12) );
  NOR2_X1 U695 ( .A1(n617), .A2(n621), .ZN(n619) );
  XNOR2_X1 U696 ( .A(G128), .B(KEYINPUT29), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n619), .B(n618), .ZN(G30) );
  XOR2_X1 U698 ( .A(G143), .B(n620), .Z(G45) );
  NOR2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U700 ( .A(G146), .B(n623), .Z(G48) );
  NAND2_X1 U701 ( .A1(n626), .A2(n624), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(G113), .ZN(G15) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(G116), .ZN(G18) );
  XOR2_X1 U705 ( .A(KEYINPUT111), .B(KEYINPUT37), .Z(n631) );
  XNOR2_X1 U706 ( .A(G125), .B(n629), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(G27) );
  XOR2_X1 U708 ( .A(G140), .B(n632), .Z(G42) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT80), .ZN(n636) );
  AND2_X1 U710 ( .A1(n710), .A2(n634), .ZN(n635) );
  OR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n669), .A2(n647), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n648), .B(KEYINPUT114), .ZN(n665) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT50), .ZN(n658) );
  NOR2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(n654), .Z(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U723 ( .A(KEYINPUT51), .B(n661), .Z(n663) );
  NAND2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U726 ( .A(n668), .B(KEYINPUT115), .ZN(n671) );
  NAND2_X1 U727 ( .A1(n669), .A2(n662), .ZN(n670) );
  XNOR2_X1 U728 ( .A(KEYINPUT53), .B(n672), .ZN(G75) );
  NAND2_X1 U729 ( .A1(n692), .A2(G469), .ZN(n673) );
  XOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n676) );
  XNOR2_X1 U731 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n675) );
  XNOR2_X1 U732 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n696), .A2(n679), .ZN(G54) );
  XNOR2_X1 U735 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT59), .ZN(n681) );
  XOR2_X1 U737 ( .A(n681), .B(KEYINPUT84), .Z(n684) );
  XNOR2_X1 U738 ( .A(n682), .B(KEYINPUT66), .ZN(n683) );
  XNOR2_X1 U739 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U740 ( .A(KEYINPUT60), .B(n686), .ZN(G60) );
  XNOR2_X1 U741 ( .A(n687), .B(KEYINPUT122), .ZN(n689) );
  NAND2_X1 U742 ( .A1(G478), .A2(n692), .ZN(n688) );
  XNOR2_X1 U743 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U744 ( .A1(n696), .A2(n690), .ZN(G63) );
  XOR2_X1 U745 ( .A(n691), .B(KEYINPUT123), .Z(n694) );
  NAND2_X1 U746 ( .A1(n692), .A2(G217), .ZN(n693) );
  XNOR2_X1 U747 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U748 ( .A1(n696), .A2(n695), .ZN(G66) );
  NAND2_X1 U749 ( .A1(G953), .A2(G224), .ZN(n697) );
  XNOR2_X1 U750 ( .A(KEYINPUT61), .B(n697), .ZN(n698) );
  NAND2_X1 U751 ( .A1(n698), .A2(G898), .ZN(n699) );
  NAND2_X1 U752 ( .A1(n700), .A2(n699), .ZN(n705) );
  XOR2_X1 U753 ( .A(n701), .B(G110), .Z(n703) );
  NOR2_X1 U754 ( .A1(G898), .A2(n711), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(KEYINPUT124), .B(n706), .ZN(G69) );
  XNOR2_X1 U758 ( .A(KEYINPUT125), .B(n707), .ZN(n709) );
  XOR2_X1 U759 ( .A(n709), .B(n708), .Z(n714) );
  XNOR2_X1 U760 ( .A(n714), .B(n710), .ZN(n712) );
  NAND2_X1 U761 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n713), .B(KEYINPUT126), .ZN(n718) );
  XNOR2_X1 U763 ( .A(G227), .B(n714), .ZN(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(G900), .ZN(n716) );
  NAND2_X1 U765 ( .A1(G953), .A2(n716), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n718), .A2(n717), .ZN(G72) );
  XNOR2_X1 U767 ( .A(G134), .B(n719), .ZN(n720) );
  XNOR2_X1 U768 ( .A(n720), .B(KEYINPUT112), .ZN(G36) );
  XOR2_X1 U769 ( .A(n721), .B(G122), .Z(G24) );
  XNOR2_X1 U770 ( .A(n722), .B(G119), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT127), .ZN(G21) );
  XOR2_X1 U772 ( .A(G131), .B(n724), .Z(G33) );
  XOR2_X1 U773 ( .A(n725), .B(G137), .Z(G39) );
endmodule

