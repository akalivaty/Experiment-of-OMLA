//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G113), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT69), .A2(G116), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(G119), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n191), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT0), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n204), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(KEYINPUT0), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT70), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G134), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n225), .A3(new_n230), .A4(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n211), .B2(new_n212), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT0), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n218), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n215), .A2(new_n241), .A3(G128), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n246), .A3(KEYINPUT1), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n245), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n215), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n243), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n226), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n223), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(G131), .C1(KEYINPUT65), .C2(new_n223), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n227), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n203), .B(new_n240), .C1(new_n258), .C2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n232), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n236), .A2(new_n238), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n258), .A2(new_n266), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n202), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n244), .A2(KEYINPUT66), .B1(new_n248), .B2(new_n250), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT68), .B(new_n215), .C1(new_n274), .C2(new_n247), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n256), .B1(new_n252), .B2(new_n253), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n242), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n265), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n203), .A4(new_n240), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n269), .A2(new_n273), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G237), .ZN(new_n281));
  INV_X1    g095(.A(G953), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(G210), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n283), .B(KEYINPUT27), .Z(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G101), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT30), .B(new_n240), .C1(new_n258), .C2(new_n266), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n214), .A2(new_n217), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n277), .A2(new_n265), .B1(new_n232), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(new_n202), .C1(new_n291), .C2(KEYINPUT30), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n286), .A3(new_n267), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n269), .A2(new_n279), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n203), .B1(new_n278), .B2(new_n240), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(KEYINPUT29), .A3(new_n287), .A4(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n296), .A2(new_n297), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G472), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n292), .A2(new_n287), .A3(new_n267), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT31), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n280), .A2(new_n286), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n292), .A2(new_n309), .A3(new_n287), .A4(new_n267), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G472), .A2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(KEYINPUT32), .A3(new_n312), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n305), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(G217), .B1(new_n318), .B2(G902), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n319), .B(KEYINPUT72), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  INV_X1    g138(.A(G221), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n325), .A2(new_n318), .A3(G953), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n324), .B(new_n326), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(G146), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n335), .A3(G146), .A4(new_n332), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n330), .A2(new_n332), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n334), .B(new_n336), .C1(G146), .C2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT67), .B(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT23), .B1(new_n216), .B2(G119), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n216), .A2(G119), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n339), .B2(G119), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT24), .B(G110), .Z(new_n346));
  AOI22_X1  g160(.A1(new_n344), .A2(G110), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n329), .A2(new_n208), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n344), .A2(G110), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n345), .A2(new_n346), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n333), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n349), .B1(new_n348), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n328), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n327), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n323), .B1(new_n359), .B2(new_n297), .ZN(new_n360));
  AOI211_X1 g174(.A(G902), .B(new_n322), .C1(new_n356), .C2(new_n358), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n321), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n319), .A2(new_n297), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n317), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(G110), .B(G140), .ZN(new_n371));
  INV_X1    g185(.A(G227), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G953), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n371), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n214), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT77), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n380), .A2(KEYINPUT77), .A3(KEYINPUT3), .A4(G104), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n386), .A3(G101), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(G101), .A3(new_n387), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n380), .A2(KEYINPUT77), .A3(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n382), .B1(new_n380), .B2(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT78), .B(G101), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n389), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n376), .B1(new_n379), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n218), .A2(new_n239), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n394), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n388), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n398), .A2(new_n401), .A3(KEYINPUT79), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n380), .A2(G104), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n384), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n393), .A2(new_n394), .B1(G101), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n277), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n242), .A2(KEYINPUT80), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n244), .A2(G128), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n253), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n242), .A2(KEYINPUT80), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n397), .A2(new_n402), .B1(new_n407), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n375), .B1(new_n415), .B2(new_n232), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n417), .A3(new_n232), .ZN(new_n418));
  INV_X1    g232(.A(new_n406), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT10), .B1(new_n258), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT79), .B1(new_n398), .B2(new_n401), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n396), .A2(new_n376), .A3(new_n218), .A4(new_n239), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT81), .B1(new_n424), .B2(new_n270), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n416), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n413), .B1(new_n277), .B2(new_n406), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT12), .B1(new_n427), .B2(new_n232), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n270), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n375), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT82), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n374), .B1(new_n424), .B2(new_n270), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n424), .A2(KEYINPUT81), .A3(new_n270), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n417), .B1(new_n415), .B2(new_n232), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  INV_X1    g253(.A(new_n430), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(new_n428), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n415), .A2(new_n232), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n374), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n434), .A2(G469), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n297), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n425), .A2(new_n418), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n375), .B1(new_n449), .B2(new_n432), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n416), .A2(new_n441), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n297), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n325), .B1(new_n455), .B2(new_n297), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n329), .B(new_n208), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n281), .A2(new_n282), .A3(G214), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n206), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n281), .A2(new_n282), .A3(G143), .A4(G214), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT18), .A2(G131), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT89), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT90), .B1(new_n464), .B2(new_n466), .ZN(new_n470));
  OAI221_X1 g284(.A(new_n460), .B1(new_n464), .B2(new_n465), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n383), .ZN(new_n473));
  AOI21_X1  g287(.A(G146), .B1(new_n330), .B2(new_n332), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(KEYINPUT73), .B2(new_n333), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(new_n263), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n463), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(KEYINPUT17), .A3(G131), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n475), .A2(new_n480), .A3(new_n481), .A4(new_n336), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n471), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n329), .B(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n333), .B1(new_n486), .B2(G146), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n479), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n333), .C1(new_n486), .C2(G146), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n473), .B1(new_n471), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n459), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT20), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n459), .C1(new_n484), .C2(new_n493), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n473), .B1(new_n471), .B2(new_n482), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n297), .B1(new_n484), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n495), .A2(new_n497), .B1(G475), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n339), .A2(G143), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n206), .A2(G128), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n219), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n503), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT92), .ZN(new_n510));
  AOI21_X1  g324(.A(G134), .B1(new_n510), .B2(new_n504), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n194), .A2(G122), .A3(new_n195), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n193), .B2(G122), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(G107), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n503), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n206), .A2(KEYINPUT13), .A3(G128), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n501), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n516), .A2(new_n517), .B1(G134), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n508), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(new_n193), .B2(G122), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G107), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n515), .B(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n505), .A2(new_n219), .A3(new_n506), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(new_n511), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n455), .A2(G217), .A3(new_n282), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n523), .B2(new_n528), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n297), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n531), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n539), .B(new_n297), .C1(KEYINPUT15), .C2(new_n535), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n500), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G952), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(G953), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n318), .B2(new_n281), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI211_X1 g359(.A(new_n297), .B(new_n282), .C1(G234), .C2(G237), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G214), .B1(G237), .B2(G902), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n331), .B(new_n242), .C1(new_n275), .C2(new_n276), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n271), .A2(G125), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n282), .A2(G224), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n551), .A2(KEYINPUT7), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n555));
  AOI22_X1  g369(.A1(KEYINPUT86), .A2(new_n555), .B1(new_n282), .B2(G224), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(KEYINPUT86), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n242), .A2(new_n331), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n255), .B2(new_n257), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n290), .A2(new_n331), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n196), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n198), .A2(KEYINPUT5), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(new_n187), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n406), .A2(new_n565), .A3(new_n201), .ZN(new_n566));
  XNOR2_X1  g380(.A(G110), .B(G122), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n399), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n568));
  INV_X1    g382(.A(new_n201), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n388), .B1(new_n569), .B2(new_n199), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n567), .B(KEYINPUT8), .ZN(new_n572));
  INV_X1    g386(.A(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n406), .B1(new_n201), .B2(new_n565), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n554), .A2(new_n561), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n297), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n553), .B(KEYINPUT84), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n559), .B2(new_n560), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n551), .A2(new_n552), .A3(new_n578), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n567), .B(KEYINPUT83), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n571), .A2(KEYINPUT6), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n586));
  INV_X1    g400(.A(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n202), .A2(new_n400), .A3(new_n388), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n566), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n582), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT85), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT85), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n582), .B(new_n592), .C1(new_n585), .C2(new_n589), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n577), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G210), .B1(G237), .B2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT87), .Z(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT88), .Z(new_n597));
  OR2_X1    g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n577), .B(new_n596), .C1(new_n591), .C2(new_n593), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n549), .A2(new_n550), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n458), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n370), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(new_n394), .Z(G3));
  INV_X1    g419(.A(G472), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n311), .B2(new_n297), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n313), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n366), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n458), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n596), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n591), .A2(new_n593), .ZN(new_n613));
  INV_X1    g427(.A(new_n577), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n550), .B1(new_n615), .B2(new_n599), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT94), .ZN(new_n617));
  INV_X1    g431(.A(new_n548), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT33), .B1(new_n532), .B2(new_n533), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n538), .A2(new_n620), .A3(new_n531), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n535), .A2(G902), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT95), .B(G478), .Z(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n622), .A2(new_n623), .B1(new_n534), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n500), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n550), .C1(new_n615), .C2(new_n599), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n617), .A2(new_n618), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n611), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n540), .A2(new_n537), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n499), .A2(G475), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n499), .A2(KEYINPUT96), .A3(G475), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n495), .A2(new_n497), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n635), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(new_n617), .A3(new_n618), .A4(new_n629), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT97), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n611), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n354), .A2(new_n355), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n328), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n650), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n364), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n362), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n609), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n602), .A2(new_n657), .A3(new_n457), .A4(new_n453), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT37), .B(G110), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n546), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n544), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n495), .B2(new_n497), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n634), .A2(new_n638), .A3(new_n666), .A4(new_n639), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n617), .A2(new_n629), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT100), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n294), .B2(new_n295), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n606), .B1(new_n670), .B2(new_n303), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n311), .A2(KEYINPUT32), .A3(new_n312), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n656), .B1(new_n673), .B2(new_n315), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n617), .A2(new_n675), .A3(new_n667), .A4(new_n629), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n669), .A2(new_n458), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n664), .B(KEYINPUT39), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n458), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n635), .A2(new_n500), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n550), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n685), .A2(new_n686), .A3(new_n655), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n286), .B1(new_n292), .B2(new_n267), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n267), .A2(new_n286), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n297), .B1(new_n689), .B2(new_n300), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n315), .A2(new_n316), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n601), .B(KEYINPUT38), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n682), .A2(new_n683), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n206), .ZN(G45));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n317), .A2(new_n453), .A3(new_n457), .A4(new_n655), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n626), .A2(new_n500), .A3(new_n665), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n617), .A2(new_n699), .A3(new_n629), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n617), .A2(new_n629), .A3(new_n699), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n458), .A2(new_n702), .A3(KEYINPUT101), .A4(new_n674), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  AOI21_X1  g519(.A(new_n442), .B1(new_n425), .B2(new_n418), .ZN(new_n706));
  OAI22_X1  g520(.A1(new_n706), .A2(new_n375), .B1(new_n441), .B2(new_n416), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n297), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n709), .A2(new_n452), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n317), .A3(new_n367), .A4(new_n457), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT102), .B1(new_n711), .B2(new_n630), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(new_n457), .A3(new_n452), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n368), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n630), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT103), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n718), .B(new_n720), .ZN(G15));
  NAND2_X1  g535(.A1(new_n645), .A2(new_n646), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT104), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n724), .B(new_n711), .C1(new_n645), .C2(new_n646), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n193), .ZN(G18));
  NAND2_X1  g541(.A1(new_n617), .A2(new_n629), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n713), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n674), .A2(new_n549), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n197), .ZN(G21));
  NAND3_X1  g547(.A1(new_n710), .A2(new_n457), .A3(new_n618), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n312), .B(KEYINPUT105), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n307), .A2(new_n310), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n301), .A2(new_n302), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n286), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n366), .A2(new_n740), .A3(new_n607), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n629), .A3(new_n617), .A4(new_n684), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT106), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n713), .A2(new_n548), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n728), .A2(new_n685), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NOR2_X1   g563(.A1(new_n740), .A2(new_n607), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n750), .A2(new_n655), .A3(new_n699), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n729), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  OAI21_X1  g567(.A(KEYINPUT107), .B1(new_n601), .B2(new_n686), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n598), .A2(new_n600), .A3(new_n755), .A4(new_n550), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n426), .A2(new_n433), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n447), .B1(new_n758), .B2(G469), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n452), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n457), .A3(new_n699), .A4(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n315), .A2(KEYINPUT108), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n315), .A2(KEYINPUT108), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n673), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n367), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT42), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n754), .A2(new_n457), .A3(new_n756), .ZN(new_n767));
  INV_X1    g581(.A(new_n760), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n368), .ZN(new_n770));
  INV_X1    g584(.A(new_n699), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n263), .ZN(G33));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n770), .A3(new_n667), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  NAND2_X1  g591(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G469), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n434), .B2(new_n444), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n448), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n452), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n456), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n679), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n754), .A2(new_n756), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n609), .A2(new_n655), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT110), .Z(new_n791));
  NAND2_X1  g605(.A1(new_n641), .A2(new_n636), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n626), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT43), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n789), .B1(new_n795), .B2(KEYINPUT44), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n788), .B(new_n796), .C1(KEYINPUT44), .C2(new_n795), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT111), .B(G137), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  NOR4_X1   g613(.A1(new_n789), .A2(new_n317), .A3(new_n367), .A4(new_n771), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n626), .A2(new_n792), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n618), .A3(new_n541), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n601), .A2(new_n550), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n610), .A3(new_n457), .A4(new_n453), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n658), .B(new_n809), .C1(new_n730), .C2(new_n731), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n748), .A3(new_n718), .A4(new_n604), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n640), .A2(new_n634), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n666), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n666), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n789), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n698), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n818), .A2(new_n819), .B1(new_n769), .B2(new_n751), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n766), .A2(new_n820), .A3(new_n773), .A4(new_n776), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n726), .A2(new_n812), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n362), .A2(new_n457), .A3(new_n654), .A4(new_n664), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n692), .A2(new_n760), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n745), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n677), .A2(new_n752), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n830), .B2(new_n704), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n729), .A2(new_n751), .B1(new_n745), .B2(new_n828), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n704), .A2(KEYINPUT114), .A3(new_n832), .A4(new_n677), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n826), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n701), .A2(new_n703), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n677), .A2(new_n752), .A3(new_n829), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(new_n841), .B2(new_n833), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n677), .A2(new_n752), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n829), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n825), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n833), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT115), .B1(new_n848), .B2(new_n826), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n836), .B(KEYINPUT52), .C1(new_n841), .C2(new_n833), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n825), .B(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n824), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(new_n826), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n822), .B1(new_n855), .B2(new_n842), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n822), .B(KEYINPUT53), .C1(new_n855), .C2(new_n842), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n822), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n867), .B2(new_n851), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n868), .B2(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n870));
  INV_X1    g684(.A(new_n710), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n871), .A2(new_n767), .A3(new_n544), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n794), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n367), .A3(new_n764), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT48), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n794), .A2(new_n545), .A3(new_n741), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n543), .B1(new_n730), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n692), .A2(new_n366), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n880), .B2(new_n627), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n873), .A2(new_n655), .A3(new_n750), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n626), .A2(new_n500), .ZN(new_n883));
  INV_X1    g697(.A(new_n876), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n693), .A2(new_n550), .A3(new_n713), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(KEYINPUT50), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT50), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OAI221_X1 g701(.A(new_n882), .B1(new_n879), .B2(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n801), .A2(new_n802), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n457), .B2(new_n871), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n876), .A2(new_n789), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n875), .B(new_n881), .C1(new_n892), .C2(KEYINPUT51), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(KEYINPUT51), .B2(new_n892), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n854), .A4(new_n858), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n861), .A2(new_n870), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n542), .A2(new_n282), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n793), .A2(new_n457), .A3(new_n550), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n366), .B(new_n899), .C1(new_n871), .C2(KEYINPUT49), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT112), .Z(new_n901));
  NOR2_X1   g715(.A1(new_n693), .A2(new_n692), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n901), .B(new_n902), .C1(KEYINPUT49), .C2(new_n871), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n898), .A2(new_n903), .ZN(G75));
  OR2_X1    g718(.A1(new_n585), .A2(new_n589), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n582), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n823), .B1(new_n867), .B2(new_n851), .ZN(new_n909));
  INV_X1    g723(.A(new_n858), .ZN(new_n910));
  OAI21_X1  g724(.A(G902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n596), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n914), .B(new_n908), .C1(new_n911), .C2(new_n597), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n282), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(new_n447), .B(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n854), .B1(new_n853), .B2(new_n858), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT54), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n707), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n911), .A2(new_n780), .A3(new_n779), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(G54));
  NOR2_X1   g741(.A1(new_n484), .A2(new_n493), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n929), .B1(new_n912), .B2(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n911), .A2(new_n928), .A3(new_n930), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n917), .A3(new_n933), .ZN(G60));
  INV_X1    g748(.A(new_n622), .ZN(new_n935));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n922), .B2(new_n923), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n918), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n861), .A2(new_n870), .A3(new_n895), .ZN(new_n941));
  INV_X1    g755(.A(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n943), .B2(new_n935), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n653), .B(new_n947), .C1(new_n909), .C2(new_n910), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n853), .B2(new_n858), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n918), .B(new_n948), .C1(new_n949), .C2(new_n359), .ZN(new_n950));
  NAND2_X1  g764(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n947), .B1(new_n909), .B2(new_n910), .ZN(new_n956));
  INV_X1    g770(.A(new_n359), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n917), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(new_n952), .A3(new_n953), .A4(new_n948), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n955), .A2(new_n959), .ZN(G66));
  NOR2_X1   g774(.A1(new_n726), .A2(new_n812), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT121), .ZN(new_n962));
  NAND2_X1  g776(.A1(G224), .A2(G953), .ZN(new_n963));
  OAI22_X1  g777(.A1(new_n962), .A2(G953), .B1(new_n547), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(G898), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n905), .B1(new_n965), .B2(G953), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  NAND4_X1  g781(.A1(new_n788), .A2(new_n367), .A3(new_n745), .A4(new_n764), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n766), .A2(new_n773), .A3(new_n776), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n845), .A2(new_n704), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n797), .A2(new_n968), .A3(new_n803), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n289), .B1(new_n291), .B2(KEYINPUT30), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n486), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n662), .B2(new_n282), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT124), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n797), .A2(new_n803), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n757), .A2(new_n541), .A3(new_n805), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n370), .A2(new_n979), .A3(new_n680), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n695), .A2(new_n970), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n983), .A2(KEYINPUT123), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(KEYINPUT123), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n978), .B(new_n982), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n282), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n975), .B(KEYINPUT122), .Z(new_n988));
  AOI21_X1  g802(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(G953), .B1(new_n372), .B2(new_n662), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G72));
  XNOR2_X1  g805(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n606), .A2(new_n297), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n992), .B(new_n993), .Z(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n962), .B2(new_n972), .ZN(new_n996));
  INV_X1    g810(.A(new_n293), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n917), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT126), .Z(new_n999));
  NOR3_X1   g813(.A1(new_n997), .A2(new_n688), .A3(new_n994), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n869), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n995), .B1(new_n986), .B2(new_n962), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n688), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(G57));
endmodule


