//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1308,
    new_n1309, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368;
  OR2_X1    g0000(.A1(KEYINPUT64), .A2(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(KEYINPUT64), .A2(G50), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n206), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n215), .A2(new_n216), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  INV_X1    g0026(.A(new_n202), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n210), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT0), .Z(new_n236));
  NOR4_X1   g0036(.A1(new_n225), .A2(new_n226), .A3(new_n233), .A4(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT69), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT73), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(KEYINPUT73), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n258), .A2(new_n230), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n231), .A2(G1), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(G68), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT11), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n258), .A2(new_n230), .A3(new_n259), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G50), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n270), .A2(new_n271), .B1(new_n231), .B2(G68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n231), .A2(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n268), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n266), .B1(new_n267), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n276), .A2(new_n267), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n261), .A2(G68), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT12), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI211_X1 g0085(.A(G226), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(G232), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT78), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT78), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT70), .B(G41), .ZN(new_n297));
  INV_X1    g0097(.A(G45), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n260), .A2(G274), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT79), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n297), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT79), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  INV_X1    g0107(.A(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(G1), .B(G13), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n304), .A2(new_n306), .B1(G238), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n295), .A2(new_n296), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n296), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n309), .B1(new_n291), .B2(new_n292), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n305), .A2(KEYINPUT79), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n303), .B(new_n300), .C1(new_n297), .C2(new_n298), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n315), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(KEYINPUT81), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT81), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(new_n315), .C1(new_n316), .C2(new_n320), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(G169), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n322), .A2(new_n324), .A3(new_n327), .A4(G169), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n316), .B2(new_n320), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n314), .A2(G179), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n282), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n248), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT74), .B(G58), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n334), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n264), .ZN(new_n338));
  INV_X1    g0138(.A(new_n261), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n263), .B1(new_n339), .B2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n258), .A2(new_n230), .A3(new_n259), .ZN(new_n342));
  INV_X1    g0142(.A(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n227), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT82), .B(G33), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n285), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT3), .ZN(new_n352));
  OR2_X1    g0152(.A1(KEYINPUT82), .A2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT82), .A2(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT83), .B1(new_n355), .B2(new_n285), .ZN(new_n356));
  AND2_X1   g0156(.A1(KEYINPUT82), .A2(G33), .ZN(new_n357));
  NOR2_X1   g0157(.A1(KEYINPUT82), .A2(G33), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT3), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT83), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n352), .A2(new_n307), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(G20), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n351), .B1(new_n363), .B2(KEYINPUT7), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n346), .B1(new_n364), .B2(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n342), .B1(new_n365), .B2(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT3), .A2(G33), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n350), .C1(new_n347), .C2(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n361), .A2(new_n367), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n349), .B1(new_n369), .B2(G20), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n345), .B1(new_n371), .B2(new_n343), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n341), .B1(new_n366), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G226), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G223), .B2(G1698), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n361), .B2(new_n359), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n307), .A2(new_n212), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n294), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n305), .B1(new_n312), .B2(G232), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G179), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(G169), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT18), .B1(new_n375), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n351), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n355), .A2(KEYINPUT83), .A3(new_n285), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n231), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(new_n349), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT16), .B(new_n345), .C1(new_n392), .C2(new_n343), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n268), .A3(new_n374), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n386), .B1(new_n394), .B2(new_n340), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT84), .ZN(new_n398));
  INV_X1    g0198(.A(G190), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n381), .A2(new_n399), .A3(new_n382), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(G200), .B1(new_n381), .B2(new_n382), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n402), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT84), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n394), .A2(new_n406), .A3(new_n340), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n394), .A2(new_n406), .A3(KEYINPUT17), .A4(new_n340), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n387), .A2(new_n397), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT8), .A2(G58), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n335), .A2(new_n269), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G20), .A2(G77), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(KEYINPUT75), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n273), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT75), .B1(new_n413), .B2(new_n414), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n268), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g0221(.A(KEYINPUT76), .B(new_n268), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n262), .A2(new_n274), .A3(new_n264), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n274), .B2(new_n339), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G244), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n302), .B1(new_n427), .B2(new_n311), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n369), .A2(G232), .A3(new_n283), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n284), .A2(new_n285), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G107), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n369), .A2(G1698), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n429), .B(new_n431), .C1(new_n432), .C2(new_n319), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n294), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G190), .ZN(new_n435));
  INV_X1    g0235(.A(G200), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(new_n434), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n294), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n305), .B1(new_n312), .B2(G244), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n384), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n434), .B2(G169), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n423), .B2(new_n425), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n369), .A2(G222), .A3(new_n283), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n430), .A2(G77), .ZN(new_n446));
  XOR2_X1   g0246(.A(KEYINPUT72), .B(G223), .Z(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n432), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n294), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n302), .B(KEYINPUT71), .C1(new_n376), .C2(new_n311), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT71), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n311), .A2(new_n376), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(new_n305), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(G179), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n273), .B2(new_n337), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(new_n268), .B1(new_n271), .B2(new_n339), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n263), .A2(G50), .A3(new_n265), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G169), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT10), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT9), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n460), .A2(new_n465), .B1(new_n454), .B2(G200), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n458), .A2(KEYINPUT9), .A3(new_n459), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n449), .A2(new_n450), .A3(new_n453), .A4(G190), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT77), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n464), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n464), .A2(new_n471), .A3(new_n467), .A4(new_n466), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n444), .B(new_n463), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n322), .A2(G200), .A3(new_n324), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n314), .A2(G190), .A3(new_n329), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n281), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR4_X1   g0278(.A1(new_n333), .A2(new_n411), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT88), .B(KEYINPUT22), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n212), .A2(G20), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n369), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(G20), .B(new_n212), .C1(new_n359), .C2(new_n361), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n231), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n347), .A2(G116), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(G20), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n480), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n231), .B(G87), .C1(new_n355), .C2(new_n285), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n483), .B1(new_n496), .B2(KEYINPUT22), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n497), .A2(KEYINPUT24), .A3(new_n493), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n268), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n260), .A2(G33), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n262), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n207), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n339), .A2(new_n207), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT25), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n499), .A2(KEYINPUT89), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT89), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT24), .B1(new_n497), .B2(new_n493), .ZN(new_n510));
  AOI21_X1  g0310(.A(G20), .B1(new_n359), .B2(new_n361), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n486), .B1(new_n511), .B2(G87), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n480), .B(new_n494), .C1(new_n512), .C2(new_n483), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n342), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n507), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n214), .A2(G1698), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G250), .B2(G1698), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n361), .B2(new_n359), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n357), .A2(new_n358), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n294), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G41), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT5), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n298), .A2(G1), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n524), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(KEYINPUT85), .B(new_n529), .C1(new_n297), .C2(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n309), .A2(G274), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n529), .B(new_n533), .C1(new_n297), .C2(KEYINPUT5), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G264), .A3(new_n309), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n523), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G169), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n384), .B2(new_n538), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n508), .A2(new_n516), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(G200), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n399), .B2(new_n538), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n514), .A3(new_n515), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n502), .A2(G87), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n359), .A2(new_n361), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n231), .A3(G68), .ZN(new_n550));
  NOR2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n212), .B1(new_n288), .B2(new_n231), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G97), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n552), .A2(new_n553), .B1(new_n273), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n342), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n416), .A2(new_n339), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n548), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n319), .A2(new_n283), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n427), .A2(G1698), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n359), .B2(new_n361), .ZN(new_n564));
  INV_X1    g0364(.A(G116), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n520), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n560), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(KEYINPUT86), .B(new_n492), .C1(new_n348), .C2(new_n563), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n294), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n529), .A2(new_n213), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n300), .A2(new_n298), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n309), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(KEYINPUT87), .B(new_n559), .C1(new_n573), .C2(new_n436), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n572), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n399), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n436), .B1(new_n569), .B2(new_n572), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n550), .A2(new_n555), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n557), .B(new_n547), .C1(new_n580), .C2(new_n342), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  OAI221_X1 g0383(.A(new_n557), .B1(new_n416), .B2(new_n503), .C1(new_n580), .C2(new_n342), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n569), .A2(G179), .A3(new_n572), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n461), .B1(new_n569), .B2(new_n572), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n342), .A2(G116), .A3(new_n261), .A4(new_n500), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n339), .A2(new_n565), .ZN(new_n591));
  AOI21_X1  g0391(.A(G20), .B1(G33), .B2(G283), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n307), .A2(G97), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(new_n593), .B1(G20), .B2(new_n565), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n268), .A2(KEYINPUT20), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT20), .B1(new_n268), .B2(new_n594), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n590), .B(new_n591), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n214), .A2(new_n283), .ZN(new_n599));
  INV_X1    g0399(.A(G264), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n359), .B2(new_n361), .ZN(new_n603));
  INV_X1    g0403(.A(G303), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n369), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n294), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n536), .A2(G270), .A3(new_n309), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n535), .A2(new_n606), .A3(G179), .A4(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n535), .A2(new_n606), .A3(new_n607), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n597), .A3(G169), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n610), .A2(new_n597), .A3(new_n613), .A4(G169), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n427), .A2(G1698), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n348), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n616), .A2(new_n427), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n620), .B(new_n283), .C1(new_n285), .C2(new_n284), .ZN(new_n621));
  OAI211_X1 g0421(.A(G250), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n622));
  NAND2_X1  g0422(.A1(G33), .A2(G283), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n309), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n536), .A2(G257), .A3(new_n309), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n535), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G169), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT4), .B1(new_n549), .B2(new_n617), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n294), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(G179), .A3(new_n535), .A4(new_n626), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(G97), .A2(G107), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT6), .B1(new_n208), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI22_X1  g0437(.A1(new_n637), .A2(new_n231), .B1(new_n274), .B2(new_n270), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n207), .B1(new_n368), .B2(new_n370), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n268), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n502), .A2(G97), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n261), .A2(G97), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n633), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n631), .A2(G190), .A3(new_n535), .A4(new_n626), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n625), .B2(new_n627), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n597), .B1(new_n610), .B2(G200), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n399), .B2(new_n610), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n615), .A2(new_n645), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n589), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n479), .A2(new_n546), .A3(new_n653), .ZN(G372));
  INV_X1    g0454(.A(new_n463), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n409), .A2(new_n410), .ZN(new_n656));
  INV_X1    g0456(.A(new_n478), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n423), .A2(new_n425), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT93), .B1(new_n658), .B2(new_n442), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n443), .A2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n656), .B1(new_n662), .B2(new_n333), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n395), .B(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n472), .A2(new_n473), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n479), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n586), .A2(new_n587), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n575), .A2(G169), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT90), .B1(new_n671), .B2(new_n585), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n584), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n645), .A2(new_n649), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n559), .B1(new_n573), .B2(new_n436), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(new_n576), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n674), .A3(new_n545), .A4(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n499), .A2(new_n507), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n540), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n615), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n675), .A2(new_n576), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n669), .B1(new_n586), .B2(new_n587), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n671), .A2(KEYINPUT90), .A3(new_n585), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n584), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n645), .A2(new_n649), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n544), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(KEYINPUT91), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n679), .A2(new_n682), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n645), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n583), .A2(new_n588), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n628), .A2(new_n632), .A3(KEYINPUT92), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT92), .B1(new_n628), .B2(new_n632), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(new_n646), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT26), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n673), .A2(new_n697), .A3(new_n698), .A4(new_n676), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n694), .A2(new_n699), .A3(new_n673), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n667), .B1(new_n668), .B2(new_n701), .ZN(G369));
  NAND3_X1  g0502(.A1(new_n260), .A2(new_n231), .A3(G13), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n680), .A2(new_n540), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n615), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n709), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n541), .A2(new_n709), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n508), .A2(new_n516), .A3(new_n708), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n541), .A2(new_n716), .A3(new_n545), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n711), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n598), .A2(new_n709), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n615), .B(new_n651), .C1(new_n598), .C2(new_n709), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n297), .ZN(new_n727));
  INV_X1    g0527(.A(new_n234), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n732), .A2(KEYINPUT95), .B1(new_n228), .B2(new_n730), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(KEYINPUT95), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  AND3_X1   g0535(.A1(new_n645), .A2(new_n649), .A3(KEYINPUT98), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT98), .B1(new_n645), .B2(new_n649), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n541), .A2(new_n615), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n545), .A3(new_n687), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n693), .A2(new_n698), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n673), .A2(new_n697), .A3(KEYINPUT26), .A4(new_n676), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n743), .A3(new_n673), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT29), .A3(new_n709), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n708), .B1(new_n691), .B2(new_n700), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n535), .A2(new_n606), .A3(new_n607), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n523), .A2(new_n537), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n572), .A4(new_n569), .ZN(new_n752));
  OAI21_X1  g0552(.A(KEYINPUT30), .B1(new_n752), .B2(new_n632), .ZN(new_n753));
  INV_X1    g0553(.A(new_n632), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n523), .A2(new_n537), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n610), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n754), .A2(new_n573), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n384), .B1(new_n625), .B2(new_n627), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n538), .A2(new_n610), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n753), .A2(new_n758), .B1(new_n761), .B2(new_n575), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT96), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n708), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n753), .A2(new_n758), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n575), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n765), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n749), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n653), .A2(new_n546), .A3(new_n709), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n766), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G330), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n748), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n735), .B1(new_n775), .B2(G1), .ZN(G364));
  NOR2_X1   g0576(.A1(new_n231), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n399), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n207), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n399), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n384), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n369), .B1(new_n783), .B2(new_n206), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n779), .B(new_n784), .C1(G87), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(G20), .A2(G179), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT100), .Z(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n399), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n436), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n787), .B1(new_n343), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n777), .A2(new_n399), .A3(new_n436), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n399), .A2(new_n436), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n789), .A2(new_n780), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n798), .B1(new_n271), .B2(new_n800), .C1(new_n336), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n790), .A2(G200), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n793), .B(new_n802), .C1(G77), .C2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT102), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT102), .ZN(new_n806));
  INV_X1    g0606(.A(G329), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n430), .B1(new_n794), .B2(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n783), .A2(new_n521), .B1(new_n785), .B2(new_n604), .ZN(new_n809));
  INV_X1    g0609(.A(new_n778), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n808), .B(new_n809), .C1(G283), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G311), .A2(new_n803), .B1(new_n791), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n801), .ZN(new_n814));
  INV_X1    g0614(.A(new_n800), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G322), .A2(new_n814), .B1(new_n815), .B2(G326), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n805), .A2(new_n806), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n230), .B1(G20), .B2(new_n461), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n722), .A2(new_n723), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n728), .A2(new_n430), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G355), .B1(new_n565), .B2(new_n728), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n251), .A2(new_n298), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n389), .A2(new_n390), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n728), .ZN(new_n829));
  INV_X1    g0629(.A(new_n229), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(G45), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n823), .A2(new_n819), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G13), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G45), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(KEYINPUT99), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(G1), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n729), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n820), .A2(new_n824), .A3(new_n834), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n724), .A2(new_n841), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n722), .A2(new_n723), .A3(new_n720), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  OAI21_X1  g0647(.A(new_n444), .B1(new_n658), .B2(new_n709), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n659), .A2(new_n661), .A3(new_n426), .A4(new_n708), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n746), .A2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n708), .B(new_n850), .C1(new_n691), .C2(new_n700), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n841), .B1(new_n855), .B2(new_n773), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n773), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n819), .A2(new_n821), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n841), .B1(G77), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n778), .A2(new_n212), .ZN(new_n861));
  INV_X1    g0661(.A(G311), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n430), .B1(new_n794), .B2(new_n862), .C1(new_n783), .C2(new_n206), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(G107), .C2(new_n786), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G294), .A2(new_n814), .B1(new_n815), .B2(G303), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT103), .B(G283), .Z(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G116), .A2(new_n803), .B1(new_n791), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G137), .A2(new_n815), .B1(new_n814), .B2(G143), .ZN(new_n870));
  INV_X1    g0670(.A(new_n803), .ZN(new_n871));
  INV_X1    g0671(.A(G150), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n871), .B2(new_n795), .C1(new_n872), .C2(new_n792), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT34), .ZN(new_n875));
  INV_X1    g0675(.A(new_n828), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n778), .A2(new_n343), .B1(new_n794), .B2(new_n877), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n783), .A2(new_n336), .B1(new_n785), .B2(new_n271), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n874), .A2(KEYINPUT34), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n869), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n860), .B1(new_n883), .B2(new_n819), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n822), .B2(new_n851), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n836), .A2(new_n260), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n345), .B1(new_n392), .B2(new_n343), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n373), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n341), .B1(new_n366), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n407), .B1(new_n890), .B2(new_n706), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n386), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n394), .A2(new_n340), .ZN(new_n894));
  INV_X1    g0694(.A(new_n386), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n706), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n898), .A3(new_n899), .A4(new_n407), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n890), .A2(new_n706), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n411), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT38), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n896), .A2(new_n898), .A3(new_n407), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n898), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n900), .A2(new_n906), .B1(new_n411), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n904), .B1(new_n908), .B2(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n770), .A2(KEYINPUT96), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n762), .A2(new_n763), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n910), .A2(KEYINPUT31), .A3(new_n708), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n768), .A2(new_n912), .A3(new_n769), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n281), .A2(new_n709), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n332), .A2(new_n657), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n330), .A3(new_n328), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n282), .B(new_n708), .C1(new_n918), .C2(new_n478), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n913), .A2(new_n920), .A3(new_n851), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n893), .A2(new_n900), .ZN(new_n924));
  INV_X1    g0724(.A(new_n902), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n664), .B2(new_n656), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT40), .B1(new_n927), .B2(new_n904), .ZN(new_n928));
  AOI22_X1  g0728(.A1(KEYINPUT40), .A2(new_n922), .B1(new_n928), .B2(new_n921), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n479), .A2(new_n913), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(G330), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n443), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n708), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n746), .B2(new_n851), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n927), .A2(new_n904), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(new_n920), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT38), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n906), .A2(new_n900), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n411), .A2(new_n907), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n927), .A2(KEYINPUT39), .A3(new_n904), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n332), .A2(new_n708), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n664), .A2(new_n897), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n479), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n667), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n887), .B1(new_n934), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n934), .ZN(new_n956));
  INV_X1    g0756(.A(new_n637), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(KEYINPUT35), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n958), .A2(G116), .A3(new_n232), .A4(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  INV_X1    g0761(.A(new_n336), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n274), .B(new_n228), .C1(new_n962), .C2(G68), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n201), .A2(new_n203), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n343), .ZN(new_n965));
  OAI211_X1 g0765(.A(G1), .B(new_n835), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n961), .A3(new_n966), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n581), .A2(new_n708), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n673), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n687), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n644), .A2(new_n708), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT98), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n688), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n645), .A2(new_n649), .A3(KEYINPUT98), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n974), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n975), .A2(new_n981), .B1(new_n697), .B2(new_n708), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n645), .B1(new_n982), .B2(new_n541), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n709), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n714), .A2(new_n718), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n982), .A2(new_n985), .A3(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT42), .B1(new_n982), .B2(new_n985), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n973), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n973), .A3(new_n989), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n982), .A2(new_n725), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n992), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n995), .A2(new_n990), .B1(new_n725), .B2(new_n982), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n729), .B(KEYINPUT41), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n975), .A2(new_n981), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n697), .A2(new_n708), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n719), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n719), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n985), .ZN(new_n1007));
  OAI211_X1 g0807(.A(KEYINPUT44), .B(new_n982), .C1(new_n1007), .C2(new_n711), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1000), .B2(new_n719), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n725), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n718), .A2(new_n724), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1014), .A2(new_n725), .A3(new_n714), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n714), .B1(new_n1014), .B2(new_n725), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n774), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1006), .A2(new_n1011), .A3(new_n725), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1013), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n997), .B1(new_n1019), .B2(new_n775), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n994), .B(new_n996), .C1(new_n1020), .C2(new_n840), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n970), .A2(new_n823), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n800), .A2(new_n862), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n785), .A2(new_n565), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n801), .A2(new_n604), .B1(new_n1024), .B2(KEYINPUT46), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(KEYINPUT46), .C2(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n783), .A2(new_n207), .B1(new_n1027), .B2(new_n794), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G97), .B2(new_n810), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G294), .A2(new_n791), .B1(new_n803), .B2(new_n867), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n876), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G159), .A2(new_n791), .B1(new_n803), .B2(new_n964), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n783), .A2(new_n343), .ZN(new_n1033));
  INV_X1    g0833(.A(G137), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n369), .B1(new_n794), .B2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n274), .A2(new_n778), .B1(new_n785), .B2(new_n336), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G143), .A2(new_n815), .B1(new_n814), .B2(G150), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1032), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n819), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n829), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n833), .B1(new_n234), .B2(new_n416), .C1(new_n1043), .C2(new_n245), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n841), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1022), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1021), .A2(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n715), .A2(new_n717), .A3(new_n823), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n825), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1051), .A2(new_n731), .B1(G107), .B2(new_n234), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n241), .A2(new_n298), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n335), .A2(new_n412), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n271), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT50), .Z(new_n1057));
  INV_X1    g0857(.A(new_n731), .ZN(new_n1058));
  AOI211_X1 g0858(.A(G45), .B(new_n1058), .C1(G68), .C2(G77), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1043), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1052), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n833), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n841), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n828), .B1(new_n871), .B2(new_n343), .C1(new_n337), .C2(new_n792), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n783), .A2(new_n416), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G77), .B2(new_n786), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n206), .B2(new_n778), .C1(new_n872), .C2(new_n794), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n271), .A2(new_n801), .B1(new_n800), .B2(new_n795), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n1064), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G317), .A2(new_n814), .B1(new_n815), .B2(G322), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n871), .B2(new_n604), .C1(new_n862), .C2(new_n792), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n782), .A2(new_n867), .B1(new_n786), .B2(G294), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT49), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n778), .A2(new_n565), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n794), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1079), .B(new_n828), .C1(G326), .C2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1069), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1063), .B1(new_n1083), .B2(new_n819), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1049), .A2(new_n840), .B1(new_n1050), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1017), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n729), .B(KEYINPUT108), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n775), .A2(new_n1049), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(G393));
  AND3_X1   g0890(.A1(new_n1006), .A2(new_n1011), .A3(new_n725), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n1012), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n840), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n369), .B(new_n779), .C1(G322), .C2(new_n1080), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n786), .A2(new_n867), .B1(new_n782), .B2(G116), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n604), .C2(new_n792), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n862), .A2(new_n801), .B1(new_n800), .B2(new_n1027), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1098));
  XNOR2_X1  g0898(.A(new_n1097), .B(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(G294), .C2(new_n803), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT111), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n872), .A2(new_n800), .B1(new_n801), .B2(new_n795), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  AOI22_X1  g0903(.A1(G68), .A2(new_n786), .B1(new_n1080), .B2(G143), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT109), .Z(new_n1105));
  NOR2_X1   g0905(.A1(new_n783), .A2(new_n274), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n876), .A2(new_n861), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n964), .A2(new_n791), .B1(new_n803), .B2(new_n1055), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1101), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT112), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n819), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n982), .A2(new_n823), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n841), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n829), .A2(new_n254), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1062), .B1(G97), .B2(new_n728), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT113), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1092), .B2(new_n1017), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1086), .B(KEYINPUT113), .C1(new_n1091), .C2(new_n1012), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1019), .A2(new_n1087), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1119), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G390));
  NAND4_X1  g0927(.A1(new_n772), .A2(new_n920), .A3(G330), .A4(new_n851), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(KEYINPUT116), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(KEYINPUT116), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n948), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n920), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n937), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n946), .A2(new_n947), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n744), .A2(new_n851), .A3(new_n709), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n936), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n916), .A2(KEYINPUT114), .A3(new_n919), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT114), .B1(new_n916), .B2(new_n919), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n394), .A2(new_n406), .A3(new_n340), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n395), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n899), .B1(new_n1146), .B2(new_n898), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n900), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n898), .B1(new_n664), .B2(new_n656), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n923), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n948), .B1(new_n1151), .B2(new_n904), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1143), .A2(new_n1144), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1144), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1131), .B(new_n1136), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n920), .B1(new_n853), .B2(new_n936), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(new_n1132), .B1(new_n946), .B2(new_n947), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1143), .A2(new_n1152), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT115), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1143), .A2(new_n1152), .A3(new_n1144), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n913), .A2(new_n920), .A3(G330), .A4(new_n851), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1155), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n840), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1114), .B1(new_n337), .B2(new_n858), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT119), .Z(new_n1167));
  OAI221_X1 g0967(.A(new_n430), .B1(new_n794), .B2(new_n521), .C1(new_n212), .C2(new_n785), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1106), .B(new_n1168), .C1(G68), .C2(new_n810), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G116), .A2(new_n814), .B1(new_n815), .B2(G283), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n803), .B1(new_n791), .B2(G107), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n1173), .A2(new_n800), .B1(new_n801), .B2(new_n877), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT120), .Z(new_n1175));
  AOI21_X1  g0975(.A(new_n430), .B1(new_n1080), .B2(G125), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n964), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n778), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G159), .B2(new_n782), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n785), .A2(new_n872), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT54), .B(G143), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n803), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n791), .A2(G137), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1172), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1167), .B1(new_n1186), .B2(new_n819), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1135), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n822), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1165), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT117), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n479), .A2(new_n1191), .A3(G330), .A4(new_n913), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n333), .A2(new_n478), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n411), .A2(new_n474), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n913), .A2(G330), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT117), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n667), .A3(new_n952), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1133), .B1(new_n773), .B2(new_n850), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1162), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n938), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1139), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n913), .A2(G330), .A3(new_n851), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1198), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1155), .B(new_n1206), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT118), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1087), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1163), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1087), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT118), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1190), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(G378));
  NAND2_X1  g1016(.A1(new_n460), .A2(new_n897), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT55), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n666), .B2(new_n463), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n472), .A2(new_n473), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1218), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1220), .A2(new_n655), .A3(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n1219), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n922), .A2(KEYINPUT40), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT40), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n939), .A2(new_n1229), .A3(new_n921), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n720), .B(new_n1227), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n913), .A2(new_n920), .A3(new_n851), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n904), .B2(new_n1151), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT38), .B1(new_n901), .B2(new_n903), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n942), .B2(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1234), .A2(new_n1229), .B1(new_n1236), .B2(new_n1233), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1232), .B1(new_n1237), .B2(G330), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n951), .B1(new_n1231), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1227), .B1(new_n929), .B2(new_n720), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n940), .A2(new_n949), .A3(new_n950), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(G330), .A3(new_n1232), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1239), .A2(new_n840), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n841), .B1(new_n964), .B2(new_n859), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n814), .A2(G128), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n782), .A2(G150), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n786), .A2(new_n1182), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n877), .A2(new_n792), .B1(new_n871), .B2(new_n1034), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G125), .C2(new_n815), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n810), .A2(G159), .ZN(new_n1255));
  AOI211_X1 g1055(.A(G33), .B(G41), .C1(new_n1080), .C2(G124), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n876), .B1(new_n871), .B2(new_n416), .C1(new_n206), .C2(new_n792), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n727), .B(new_n1033), .C1(G283), .C2(new_n1080), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n810), .A2(new_n962), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n274), .B2(new_n785), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G107), .A2(new_n814), .B1(new_n815), .B2(G116), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1258), .A2(new_n1260), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT58), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1265), .A2(KEYINPUT58), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n271), .B1(G33), .B2(G41), .C1(new_n828), .C2(new_n727), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1257), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1245), .B1(new_n1269), .B2(new_n819), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1227), .B2(new_n822), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1244), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1198), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1207), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1239), .A2(KEYINPUT57), .A3(new_n1243), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1087), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1207), .A2(new_n1273), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1272), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT122), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(KEYINPUT122), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G375));
  INV_X1    g1083(.A(new_n997), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1205), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1210), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1164), .B1(new_n1205), .B2(new_n1201), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n821), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n841), .B1(G68), .B2(new_n859), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n430), .B1(new_n794), .B2(new_n604), .C1(new_n274), .C2(new_n778), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1065), .B(new_n1290), .C1(G97), .C2(new_n786), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G283), .A2(new_n814), .B1(new_n815), .B2(G294), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(G107), .A2(new_n803), .B1(new_n791), .B2(G116), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1294), .A2(KEYINPUT123), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n1261), .B1(new_n783), .B2(new_n271), .C1(new_n801), .C2(new_n1034), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G132), .B2(new_n815), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n803), .A2(G150), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n794), .A2(new_n1173), .B1(new_n785), .B2(new_n795), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT124), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n876), .B1(new_n791), .B2(new_n1182), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1297), .A2(new_n1298), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(KEYINPUT123), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1295), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1289), .B1(new_n1304), .B2(new_n819), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1287), .B1(new_n1288), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1286), .A2(new_n1306), .ZN(G381));
  OR3_X1    g1107(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1308));
  NOR4_X1   g1108(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1215), .B(new_n1309), .C1(new_n1281), .C2(new_n1282), .ZN(G407));
  NAND2_X1  g1110(.A1(new_n707), .A2(G213), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1215), .B(new_n1312), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(G407), .A2(new_n1313), .A3(G213), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT125), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(G407), .A2(new_n1313), .A3(new_n1316), .A4(G213), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(G409));
  NAND3_X1  g1118(.A1(new_n1277), .A2(new_n1278), .A3(new_n1284), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1272), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1214), .A2(new_n1211), .A3(new_n1209), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1190), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1280), .B2(new_n1215), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  OR2_X1    g1125(.A1(new_n1285), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1285), .A2(new_n1325), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1087), .A3(new_n1210), .A4(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1328), .A2(G384), .A3(new_n1306), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G384), .B1(new_n1328), .B2(new_n1306), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1324), .A2(new_n1311), .A3(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1324), .A2(new_n1311), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1312), .A2(G2897), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1331), .B(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1333), .A2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1324), .A2(new_n1311), .A3(new_n1331), .A4(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1334), .A2(new_n1338), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n996), .A2(new_n994), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1019), .A2(new_n775), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1284), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1344), .B1(new_n1346), .B2(new_n1164), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1126), .B1(new_n1347), .B2(new_n1046), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1124), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1021), .B(new_n1047), .C1(new_n1349), .C2(new_n1119), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(G393), .B(new_n846), .ZN(new_n1351));
  AND3_X1   g1151(.A1(new_n1348), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1351), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1343), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT126), .B1(new_n1354), .B2(new_n1339), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT126), .ZN(new_n1358));
  NOR4_X1   g1158(.A1(new_n1352), .A2(new_n1353), .A3(new_n1358), .A4(KEYINPUT61), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1324), .A2(KEYINPUT63), .A3(new_n1311), .A4(new_n1331), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT63), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1332), .A2(new_n1362), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1360), .A2(new_n1338), .A3(new_n1361), .A4(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1356), .A2(new_n1364), .ZN(G405));
  XNOR2_X1  g1165(.A(new_n1354), .B(new_n1331), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(G378), .A2(new_n1280), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1367), .B1(G375), .B2(G378), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1366), .B(new_n1368), .ZN(G402));
endmodule


