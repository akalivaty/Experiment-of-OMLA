//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT84), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT84), .A3(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT83), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(KEYINPUT82), .A3(KEYINPUT15), .ZN(new_n219));
  OR3_X1    g018(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n220), .A2(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(new_n220), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n221), .A2(new_n224), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n226), .A2(new_n227), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  OAI22_X1  g027(.A1(new_n215), .A2(new_n223), .B1(new_n216), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n210), .A2(KEYINPUT85), .A3(new_n211), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT85), .B1(new_n210), .B2(new_n211), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  OAI221_X1 g036(.A(new_n237), .B1(new_n228), .B2(new_n216), .C1(new_n215), .C2(new_n223), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n231), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n241), .B(KEYINPUT13), .Z(new_n246));
  NOR2_X1   g045(.A1(new_n212), .A2(new_n229), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT11), .B(G169gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT12), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n244), .A2(new_n245), .A3(new_n256), .A4(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT64), .Z(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  INV_X1    g061(.A(G127gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(G134gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G127gat), .ZN(new_n266));
  OAI22_X1  g065(.A1(new_n262), .A2(KEYINPUT1), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G113gat), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n282), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n277), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .A3(new_n285), .A4(new_n284), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(KEYINPUT28), .A3(new_n283), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n278), .A2(new_n283), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(KEYINPUT65), .B2(KEYINPUT24), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(KEYINPUT23), .B2(new_n295), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT23), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(new_n305), .A3(new_n306), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(new_n313), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n309), .A2(new_n315), .B1(new_n323), .B2(new_n311), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n276), .B1(new_n304), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n267), .A2(new_n275), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n327), .B(new_n324), .C1(new_n294), .C2(new_n303), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n261), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT32), .ZN(new_n330));
  XOR2_X1   g129(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G15gat), .B(G43gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n293), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n291), .A2(new_n285), .A3(new_n284), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n277), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n302), .B1(new_n340), .B2(new_n292), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n327), .B1(new_n341), .B2(new_n324), .ZN(new_n342));
  INV_X1    g141(.A(new_n261), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n304), .A2(new_n276), .A3(new_n325), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT34), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT34), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n347), .A3(new_n343), .A4(new_n344), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n336), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n329), .B(KEYINPUT32), .C1(new_n332), .C2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n337), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n337), .A2(new_n351), .B1(new_n346), .B2(new_n348), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT70), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT36), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n351), .ZN(new_n356));
  INV_X1    g155(.A(new_n349), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n370), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n369), .A2(new_n374), .A3(new_n371), .A4(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384));
  INV_X1    g183(.A(G141gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(G148gat), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n383), .A2(new_n384), .B1(new_n386), .B2(KEYINPUT73), .ZN(new_n387));
  INV_X1    g186(.A(G148gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G141gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n388), .A2(G141gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n382), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n384), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(new_n381), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n387), .A2(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT74), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n400));
  OAI22_X1  g199(.A1(new_n400), .A2(new_n395), .B1(new_n389), .B2(new_n391), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT2), .B1(new_n389), .B2(new_n390), .ZN(new_n403));
  INV_X1    g202(.A(new_n381), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n384), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT3), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n380), .B1(new_n409), .B2(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT29), .B1(new_n376), .B2(new_n377), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n411), .B2(KEYINPUT3), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n364), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n378), .A2(new_n379), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT72), .B1(new_n376), .B2(new_n377), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n406), .B2(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n397), .A2(KEYINPUT74), .A3(new_n398), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n364), .B(new_n412), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n362), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n412), .B1(new_n416), .B2(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n363), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(G22gat), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT78), .B(G22gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n427), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n413), .B2(new_n421), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n428), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n426), .A2(new_n433), .B1(new_n436), .B2(new_n431), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n397), .B(new_n327), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT5), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n276), .B1(KEYINPUT3), .B2(new_n406), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n399), .B2(new_n408), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT4), .B1(new_n276), .B2(new_n397), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n406), .A2(new_n327), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n439), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n440), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n276), .A2(new_n397), .A3(KEYINPUT4), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n444), .B1(new_n406), .B2(new_n327), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n450), .B2(new_n451), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n442), .B(new_n449), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT76), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT75), .B1(new_n443), .B2(new_n445), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n442), .A4(new_n449), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n448), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G1gat), .B(G29gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT0), .ZN(new_n464));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n462), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n461), .ZN(new_n473));
  INV_X1    g272(.A(new_n448), .ZN(new_n474));
  AND4_X1   g273(.A1(new_n473), .A2(new_n474), .A3(new_n468), .A4(new_n467), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND2_X1  g278(.A1(G226gat), .A2(G233gat), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n324), .B1(new_n294), .B2(new_n303), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(KEYINPUT29), .ZN(new_n482));
  OAI211_X1 g281(.A(G226gat), .B(G233gat), .C1(new_n341), .C2(new_n324), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n380), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n380), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n482), .A2(new_n483), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n416), .ZN(new_n491));
  INV_X1    g290(.A(new_n479), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n484), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT30), .B(new_n479), .C1(new_n485), .C2(new_n486), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n437), .B1(new_n476), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n337), .A2(new_n349), .A3(new_n351), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n358), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n361), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT80), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n474), .ZN(new_n502));
  INV_X1    g301(.A(new_n469), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n470), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n462), .A2(new_n468), .A3(new_n467), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n487), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT37), .B1(new_n485), .B2(new_n486), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n508), .A3(new_n484), .ZN(new_n509));
  AOI211_X1 g308(.A(KEYINPUT38), .B(new_n479), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n501), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT38), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT37), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n491), .B2(new_n484), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n512), .B(new_n492), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n476), .A2(KEYINPUT80), .A3(new_n515), .A4(new_n487), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n492), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT38), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n442), .B1(new_n453), .B2(new_n454), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n446), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(KEYINPUT39), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n438), .A2(new_n439), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(KEYINPUT39), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n524), .A3(new_n466), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT40), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n522), .A2(new_n524), .A3(new_n527), .A4(new_n466), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n526), .A2(new_n528), .B1(new_n502), .B2(new_n467), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n437), .B1(new_n529), .B2(new_n495), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n500), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n354), .A2(new_n360), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n476), .A2(new_n495), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n437), .A2(KEYINPUT35), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n498), .ZN(new_n537));
  INV_X1    g336(.A(new_n437), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT35), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n259), .B1(new_n532), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  OR2_X1    g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(KEYINPUT87), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n548));
  NOR2_X1   g347(.A1(G57gat), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G57gat), .A2(G64gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(KEYINPUT86), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n553));
  INV_X1    g352(.A(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n549), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n547), .A2(new_n548), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(KEYINPUT9), .A3(new_n551), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(new_n544), .A3(new_n545), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n543), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT88), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(KEYINPUT91), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n212), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT92), .ZN(new_n569));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT89), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n569), .A2(new_n575), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n565), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n577), .B2(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(KEYINPUT93), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n594), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  OR2_X1    g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT94), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n596), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT95), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n598), .A2(new_n602), .A3(new_n599), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n602), .B1(new_n598), .B2(new_n599), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n593), .B(new_n595), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n606), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n239), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n229), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n615), .A2(new_n617), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n615), .A2(new_n620), .A3(new_n617), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n621), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n560), .A2(new_n561), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n610), .A2(KEYINPUT97), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n563), .B1(new_n637), .B2(new_n606), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n610), .A2(KEYINPUT97), .A3(new_n605), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n614), .A2(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n614), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n640), .A2(new_n641), .B1(new_n567), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT98), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n635), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n647), .B(new_n641), .C1(new_n616), .C2(new_n580), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n567), .A2(new_n642), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n645), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n651), .B2(new_n640), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n657), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n651), .ZN(new_n661));
  AOI211_X1 g460(.A(new_n660), .B(new_n661), .C1(new_n650), .C2(new_n651), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n590), .A2(new_n634), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n542), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n542), .A2(KEYINPUT101), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n476), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT102), .B(G1gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n495), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n670), .ZN(new_n678));
  INV_X1    g477(.A(new_n495), .ZN(new_n679));
  OAI21_X1  g478(.A(G8gat), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(G1325gat));
  INV_X1    g481(.A(G15gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n361), .A2(new_n499), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n678), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n533), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n678), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n689), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n670), .A2(new_n437), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n542), .ZN(new_n695));
  INV_X1    g494(.A(new_n476), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n589), .A2(new_n633), .A3(new_n664), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n695), .A2(G29gat), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT45), .Z(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n361), .A2(new_n496), .A3(new_n499), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n519), .B2(new_n530), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n535), .A2(new_n534), .ZN(new_n704));
  AOI22_X1  g503(.A1(new_n704), .A2(new_n533), .B1(new_n539), .B2(KEYINPUT35), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n701), .B(new_n634), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n590), .A2(KEYINPUT104), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n590), .A2(KEYINPUT104), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n259), .A3(new_n664), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n633), .B1(new_n532), .B2(new_n541), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n714), .B2(new_n701), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT105), .B(new_n634), .C1(new_n703), .C2(new_n705), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n709), .B(new_n713), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n696), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n700), .A2(KEYINPUT107), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1328gat));
  NOR4_X1   g523(.A1(new_n695), .A2(G36gat), .A3(new_n679), .A4(new_n698), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n718), .B2(new_n679), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1329gat));
  NOR2_X1   g529(.A1(new_n695), .A2(new_n698), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n732), .A3(new_n533), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT110), .B1(new_n718), .B2(new_n685), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n718), .A2(KEYINPUT110), .A3(new_n685), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT47), .B(new_n733), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G43gat), .B1(new_n718), .B2(new_n685), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n738), .B2(new_n733), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT109), .B(KEYINPUT47), .C1(new_n738), .C2(new_n733), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(G1330gat));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  OAI21_X1  g543(.A(G50gat), .B1(new_n718), .B2(new_n538), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n695), .A2(G50gat), .A3(new_n538), .A4(new_n698), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n744), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n708), .B1(new_n714), .B2(KEYINPUT105), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n706), .A2(new_n707), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n437), .A3(new_n709), .A4(new_n713), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n746), .B1(new_n755), .B2(G50gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(KEYINPUT112), .A3(new_n749), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  AND4_X1   g557(.A1(new_n758), .A2(new_n745), .A3(KEYINPUT48), .A4(new_n747), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n756), .B2(KEYINPUT48), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n751), .A2(new_n757), .B1(new_n759), .B2(new_n760), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n532), .A2(new_n541), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n662), .B1(new_n654), .B2(new_n658), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n590), .A2(new_n258), .A3(new_n634), .A4(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n476), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g566(.A1(new_n765), .A2(new_n495), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n765), .A2(new_n684), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n687), .A2(G71gat), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n773), .A2(G71gat), .B1(new_n765), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n437), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  INV_X1    g577(.A(new_n714), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n589), .A2(new_n258), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n779), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n763), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(G85gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n787), .A3(new_n476), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n754), .A2(new_n664), .A3(new_n709), .A4(new_n781), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n696), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1336gat));
  NOR2_X1   g590(.A1(new_n679), .A2(G92gat), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT114), .B1(new_n789), .B2(new_n679), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n679), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n786), .A2(new_n792), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n789), .B2(new_n679), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n789), .B2(new_n685), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n784), .A2(new_n785), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n533), .A2(new_n664), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n805), .A2(G99gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(G1338gat));
  XNOR2_X1  g606(.A(KEYINPUT115), .B(G106gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n789), .B2(new_n538), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n538), .A2(new_n763), .A3(G106gat), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT116), .Z(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n804), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n809), .B(new_n814), .C1(new_n804), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1339gat));
  NAND2_X1  g615(.A1(new_n665), .A2(new_n259), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n646), .A2(new_n652), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n660), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT118), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n823), .A3(new_n660), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n819), .B1(new_n650), .B2(new_n651), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n650), .A2(new_n651), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n825), .B(new_n829), .C1(new_n651), .C2(new_n650), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n822), .A2(new_n824), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n634), .B1(new_n831), .B2(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n828), .A2(new_n830), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n820), .A2(new_n823), .A3(new_n660), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n823), .B1(new_n820), .B2(new_n660), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(KEYINPUT55), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n663), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n231), .A2(new_n247), .A3(new_n246), .ZN(new_n839));
  INV_X1    g638(.A(new_n234), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n239), .A2(new_n840), .A3(new_n232), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n241), .B1(new_n841), .B2(new_n230), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n240), .A2(KEYINPUT119), .A3(new_n241), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n253), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n257), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n838), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n664), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT120), .B1(new_n763), .B2(new_n847), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n259), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n662), .B1(new_n831), .B2(KEYINPUT55), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n858), .B2(new_n634), .ZN(new_n859));
  INV_X1    g658(.A(new_n712), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n818), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n696), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n537), .A2(new_n538), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n495), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n258), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n832), .A2(new_n837), .A3(new_n847), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n855), .A2(new_n854), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n258), .A3(new_n663), .A4(new_n836), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n852), .A3(new_n851), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n871), .B2(new_n633), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n817), .B1(new_n872), .B2(new_n712), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n538), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n696), .A2(new_n495), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n687), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n259), .A2(new_n270), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n867), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  AOI21_X1  g678(.A(G120gat), .B1(new_n866), .B2(new_n664), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n763), .A2(new_n268), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(G1341gat));
  INV_X1    g681(.A(new_n877), .ZN(new_n883));
  OAI21_X1  g682(.A(G127gat), .B1(new_n883), .B2(new_n860), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n263), .A3(new_n589), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1342gat));
  OAI21_X1  g685(.A(G134gat), .B1(new_n883), .B2(new_n633), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n634), .A2(new_n265), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n865), .A2(KEYINPUT56), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT56), .B1(new_n865), .B2(new_n888), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(G1343gat));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n861), .B2(new_n696), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n893), .A3(new_n476), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n684), .A2(new_n538), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n679), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n892), .A2(new_n894), .A3(new_n258), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n385), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n684), .A2(new_n876), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n259), .A2(new_n385), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n538), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n848), .A2(new_n664), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n634), .B1(new_n870), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n590), .B1(new_n906), .B2(new_n868), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n818), .B1(new_n907), .B2(KEYINPUT121), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n873), .B2(new_n437), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n900), .B(new_n901), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n899), .A2(KEYINPUT58), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n763), .A2(G148gat), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n892), .A2(new_n894), .A3(new_n897), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n847), .B1(new_n838), .B2(KEYINPUT124), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n832), .B2(new_n837), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n906), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n817), .B1(new_n925), .B2(new_n589), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n926), .B2(new_n437), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n861), .A2(new_n902), .A3(new_n538), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n664), .B(new_n900), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n921), .B1(new_n929), .B2(G148gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n921), .A2(G148gat), .ZN(new_n931));
  INV_X1    g730(.A(new_n900), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n909), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n903), .ZN(new_n934));
  INV_X1    g733(.A(new_n911), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n936), .B2(new_n664), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n920), .B1(new_n930), .B2(new_n937), .ZN(G1345gat));
  OAI21_X1  g737(.A(new_n900), .B1(new_n910), .B2(new_n911), .ZN(new_n939));
  OAI21_X1  g738(.A(G155gat), .B1(new_n939), .B2(new_n860), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n892), .A2(new_n894), .A3(new_n897), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n590), .A2(G155gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1346gat));
  NAND3_X1  g742(.A1(new_n936), .A2(G162gat), .A3(new_n634), .ZN(new_n944));
  INV_X1    g743(.A(G162gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n941), .B2(new_n633), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n944), .A2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n679), .A2(new_n476), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n863), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n873), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n258), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n874), .A2(new_n687), .A3(new_n949), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n259), .A2(new_n312), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(G1348gat));
  AOI21_X1  g755(.A(G176gat), .B1(new_n952), .B2(new_n664), .ZN(new_n957));
  INV_X1    g756(.A(new_n874), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n805), .A2(new_n313), .A3(new_n949), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(G1349gat));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n533), .A3(new_n948), .ZN(new_n961));
  OAI21_X1  g760(.A(G183gat), .B1(new_n961), .B2(new_n860), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n589), .A2(new_n287), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n962), .B(new_n963), .C1(new_n951), .C2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n278), .B1(new_n954), .B2(new_n712), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n951), .A2(new_n964), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT60), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n952), .A2(new_n283), .A3(new_n634), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n634), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(G190gat), .ZN(new_n973));
  AOI211_X1 g772(.A(KEYINPUT61), .B(new_n283), .C1(new_n954), .C2(new_n634), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n895), .A2(new_n948), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n861), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n873), .A2(KEYINPUT125), .A3(new_n895), .A4(new_n948), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(G197gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n980), .A2(new_n981), .A3(new_n258), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n684), .A2(new_n949), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n633), .B1(new_n855), .B2(new_n854), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n857), .A2(new_n985), .A3(KEYINPUT124), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n924), .A2(new_n848), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n870), .A2(new_n905), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n633), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n818), .B1(new_n990), .B2(new_n590), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n902), .B1(new_n991), .B2(new_n538), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n873), .A2(KEYINPUT57), .A3(new_n437), .ZN(new_n993));
  AOI211_X1 g792(.A(new_n259), .B(new_n984), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n995));
  OAI21_X1  g794(.A(G197gat), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n984), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(new_n995), .A3(new_n258), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n982), .B1(new_n996), .B2(new_n998), .ZN(G1352gat));
  NOR4_X1   g798(.A1(new_n861), .A2(G204gat), .A3(new_n763), .A4(new_n977), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT62), .ZN(new_n1001));
  AOI211_X1 g800(.A(new_n763), .B(new_n984), .C1(new_n992), .C2(new_n993), .ZN(new_n1002));
  INV_X1    g801(.A(G204gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G1353gat));
  NAND3_X1  g803(.A1(new_n980), .A2(new_n366), .A3(new_n589), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT63), .ZN(new_n1006));
  AOI211_X1 g805(.A(new_n1006), .B(new_n366), .C1(new_n997), .C2(new_n589), .ZN(new_n1007));
  OAI211_X1 g806(.A(new_n589), .B(new_n983), .C1(new_n927), .C2(new_n928), .ZN(new_n1008));
  AOI21_X1  g807(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1005), .B1(new_n1007), .B2(new_n1009), .ZN(G1354gat));
  NAND3_X1  g809(.A1(new_n978), .A2(new_n979), .A3(new_n634), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(new_n367), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1011), .A2(new_n1014), .A3(new_n367), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n633), .A2(new_n367), .ZN(new_n1016));
  AOI22_X1  g815(.A1(new_n1013), .A2(new_n1015), .B1(new_n997), .B2(new_n1016), .ZN(G1355gat));
endmodule


