//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G169gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G197gat), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G197gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT12), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT12), .B1(new_n206), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G22gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G15gat), .ZN(new_n215));
  INV_X1    g014(.A(G15gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G22gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n215), .A3(new_n217), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT92), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n223), .A2(G8gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n220), .B(new_n222), .C1(KEYINPUT91), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G8gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(KEYINPUT91), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT91), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n221), .A2(new_n215), .A3(new_n217), .A4(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n227), .A2(new_n228), .A3(new_n223), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G29gat), .ZN(new_n233));
  INV_X1    g032(.A(G36gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT14), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT14), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G29gat), .B2(G36gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(G29gat), .A2(G36gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT15), .ZN(new_n240));
  INV_X1    g039(.A(G43gat), .ZN(new_n241));
  INV_X1    g040(.A(G50gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G43gat), .A2(G50gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n240), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n240), .A3(new_n244), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT89), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n243), .A2(new_n249), .A3(new_n240), .A4(new_n244), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n244), .ZN(new_n252));
  NOR2_X1   g051(.A1(G43gat), .A2(G50gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT15), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n238), .A2(KEYINPUT90), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(G29gat), .A3(G36gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n258), .A3(new_n237), .A4(new_n235), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n246), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n232), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G229gat), .A2(G233gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n223), .B1(G8gat), .B2(new_n225), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n235), .A2(new_n237), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n245), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n258), .A3(new_n248), .A4(new_n250), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT17), .A3(new_n246), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT93), .A4(new_n271), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n262), .B(KEYINPUT96), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT13), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n226), .A2(new_n231), .B1(new_n270), .B2(new_n246), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT97), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n226), .A2(new_n246), .A3(new_n270), .A4(new_n231), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n276), .A2(KEYINPUT18), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n213), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT18), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n276), .B2(KEYINPUT94), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n291), .B(new_n263), .C1(new_n274), .C2(new_n275), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n286), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI221_X1 g093(.A(new_n286), .B1(new_n287), .B2(new_n213), .C1(new_n290), .C2(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(G218gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT77), .B1(new_n307), .B2(G141gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(G148gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n308), .B(new_n311), .C1(new_n310), .C2(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n316), .B2(KEYINPUT2), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n307), .A2(G141gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n310), .A2(G148gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n316), .A2(new_n313), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n306), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n312), .A2(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n305), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT29), .B1(new_n327), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n326), .B(new_n331), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT85), .B(G22gat), .Z(new_n337));
  OAI21_X1  g136(.A(new_n326), .B1(new_n327), .B2(new_n334), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n335), .A2(new_n305), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(new_n242), .ZN(new_n343));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n340), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(G22gat), .ZN(new_n350));
  AOI211_X1 g149(.A(KEYINPUT86), .B(new_n214), .C1(new_n336), .C2(new_n340), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n337), .B1(new_n336), .B2(new_n340), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n346), .B1(new_n341), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G113gat), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n359), .A2(G120gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(G120gat), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT1), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  INV_X1    g163(.A(G134gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G127gat), .ZN(new_n366));
  INV_X1    g165(.A(G127gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G134gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT67), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT67), .B1(new_n365), .B2(G127gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n364), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT67), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n366), .B2(new_n368), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n375), .A2(KEYINPUT68), .A3(new_n371), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n363), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT69), .B(G113gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G120gat), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n360), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n327), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT68), .B1(new_n375), .B2(new_n371), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n372), .B(new_n364), .C1(new_n378), .C2(new_n374), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n362), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n388), .A2(new_n325), .A3(new_n383), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n358), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n327), .A3(new_n384), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n325), .B1(new_n388), .B2(new_n383), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n357), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n384), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT78), .B1(new_n327), .B2(new_n328), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n327), .A2(new_n334), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n325), .A2(new_n401), .A3(KEYINPUT3), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n389), .A2(new_n404), .ZN(new_n405));
  NOR4_X1   g204(.A1(new_n388), .A2(new_n325), .A3(new_n383), .A4(KEYINPUT4), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n403), .B(new_n357), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n391), .A2(new_n397), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n388), .A2(new_n383), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n404), .A3(new_n327), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n412), .A2(new_n396), .A3(new_n357), .A4(new_n403), .ZN(new_n413));
  XNOR2_X1  g212(.A(G57gat), .B(G85gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT82), .B1(new_n408), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n391), .A2(new_n397), .A3(new_n407), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n413), .ZN(new_n422));
  INV_X1    g221(.A(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n427), .A3(new_n413), .A4(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n426), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n425), .A2(new_n426), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n305), .B(KEYINPUT74), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(G169gat), .A2(G176gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n442), .B1(new_n449), .B2(new_n441), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n440), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n449), .A3(new_n441), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT25), .B(new_n435), .C1(new_n438), .C2(new_n439), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n451), .A2(KEYINPUT25), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G176gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n207), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT26), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n434), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n436), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT66), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT66), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT27), .B(G183gat), .ZN(new_n464));
  INV_X1    g263(.A(G190gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(KEYINPUT28), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT28), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n462), .A2(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n456), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n433), .B1(new_n470), .B2(new_n306), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n432), .B1(new_n456), .B2(new_n469), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n431), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n454), .ZN(new_n474));
  INV_X1    g273(.A(new_n439), .ZN(new_n475));
  NOR3_X1   g274(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n434), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT64), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n478), .A2(new_n452), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n479), .A2(new_n446), .B1(new_n442), .B2(new_n441), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n449), .A2(new_n441), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT65), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n474), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n461), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT66), .ZN(new_n489));
  INV_X1    g288(.A(new_n468), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n466), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n433), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n456), .B2(new_n469), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n305), .C1(new_n493), .C2(new_n433), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT75), .B(G8gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n494), .A4(new_n499), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n306), .B1(new_n485), .B2(new_n491), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n472), .B1(new_n505), .B2(new_n432), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n494), .B(new_n499), .C1(new_n506), .C2(new_n333), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT76), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n473), .A2(new_n509), .A3(new_n494), .A4(new_n499), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n503), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT83), .B1(new_n430), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n413), .A2(new_n418), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n427), .B1(new_n514), .B2(new_n421), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n418), .B1(new_n421), .B2(new_n413), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n426), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n429), .A2(new_n424), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n512), .A4(KEYINPUT83), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n356), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n470), .B(new_n410), .ZN(new_n522));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT32), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  XOR2_X1   g325(.A(G71gat), .B(G99gat), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT70), .ZN(new_n528));
  XOR2_X1   g327(.A(G15gat), .B(G43gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n524), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  OAI221_X1 g331(.A(KEYINPUT32), .B1(new_n525), .B2(new_n530), .C1(new_n522), .C2(new_n523), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n522), .A2(KEYINPUT72), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n522), .A2(KEYINPUT72), .B1(G227gat), .B2(G233gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT34), .B1(G227gat), .B2(G233gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n522), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n522), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n532), .A2(new_n534), .B1(new_n540), .B2(new_n545), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(KEYINPUT36), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT36), .B1(new_n547), .B2(new_n548), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n517), .A2(new_n518), .A3(new_n512), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT83), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n355), .B1(new_n556), .B2(new_n519), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n549), .A2(new_n550), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n494), .B(new_n560), .C1(new_n506), .C2(new_n333), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n500), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n473), .B2(new_n494), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT38), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n560), .B1(new_n506), .B2(new_n431), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n305), .B1(new_n471), .B2(new_n472), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n561), .A3(new_n568), .A4(new_n500), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n564), .A2(new_n511), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT6), .B1(new_n420), .B2(new_n424), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n516), .B1(new_n426), .B2(new_n428), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n511), .A2(new_n504), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n502), .A3(new_n501), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n393), .A2(new_n394), .A3(new_n357), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n401), .A2(new_n329), .B1(new_n377), .B2(new_n384), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n399), .A2(new_n400), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n409), .A2(new_n411), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(KEYINPUT39), .B(new_n576), .C1(new_n579), .C2(new_n357), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n412), .A2(new_n403), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n358), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n580), .A2(new_n583), .A3(KEYINPUT40), .A4(new_n418), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT88), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n357), .B1(new_n412), .B2(new_n403), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n423), .B1(new_n587), .B2(new_n582), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n588), .A2(KEYINPUT88), .A3(new_n580), .A4(KEYINPUT40), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT40), .B1(new_n588), .B2(new_n580), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n516), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n593), .A3(new_n355), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n552), .A2(new_n559), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n547), .A2(new_n355), .A3(new_n548), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n519), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n547), .A2(new_n548), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n599), .A2(KEYINPUT35), .A3(new_n356), .ZN(new_n600));
  INV_X1    g399(.A(new_n554), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n297), .B1(new_n595), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT102), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  OR2_X1    g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(KEYINPUT101), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  INV_X1    g412(.A(G92gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT101), .B1(new_n610), .B2(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n609), .A3(new_n612), .A4(new_n615), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n267), .A2(new_n271), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n620), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n622), .A2(new_n260), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n607), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(new_n365), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n315), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n607), .A3(new_n624), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n626), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n621), .A2(KEYINPUT103), .A3(new_n624), .A4(new_n607), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G57gat), .B(G64gat), .Z(new_n644));
  NAND2_X1  g443(.A1(G71gat), .A2(G78gat), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT9), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(G71gat), .A2(G78gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(new_n645), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n644), .B(new_n647), .C1(new_n650), .C2(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n647), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n645), .A2(new_n649), .B1(new_n647), .B2(KEYINPUT98), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n232), .B1(KEYINPUT21), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT99), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(KEYINPUT21), .ZN(new_n658));
  XOR2_X1   g457(.A(G127gat), .B(G155gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  NAND2_X1  g463(.A1(G231gat), .A2(G233gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G183gat), .B(G211gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n662), .A2(new_n663), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n662), .B2(new_n663), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(G230gat), .ZN(new_n673));
  INV_X1    g472(.A(G233gat), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n622), .A2(new_n655), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n618), .A2(new_n651), .A3(new_n620), .A4(new_n654), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n655), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n676), .A2(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n675), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G120gat), .B(G148gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G176gat), .ZN(new_n687));
  INV_X1    g486(.A(G204gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n682), .A2(new_n684), .A3(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n643), .A2(new_n672), .A3(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n604), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n430), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g500(.A(KEYINPUT16), .B(G8gat), .Z(new_n702));
  NAND3_X1  g501(.A1(new_n695), .A2(new_n575), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n695), .A2(new_n575), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G8gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(G1325gat));
  AND2_X1   g508(.A1(new_n547), .A2(new_n548), .ZN(new_n710));
  AOI21_X1  g509(.A(G15gat), .B1(new_n695), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n558), .A2(G15gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT106), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n711), .B1(new_n695), .B2(new_n713), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n356), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NAND2_X1  g516(.A1(new_n595), .A2(new_n603), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n642), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n573), .A2(new_n593), .A3(new_n355), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n557), .A2(new_n722), .A3(new_n558), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n597), .A2(KEYINPUT35), .B1(new_n601), .B2(new_n600), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n643), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n719), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n672), .B(KEYINPUT108), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(new_n297), .A3(new_n693), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n721), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n699), .ZN(new_n731));
  OAI21_X1  g530(.A(G29gat), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n693), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n643), .A2(new_n672), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT107), .Z(new_n735));
  NAND4_X1  g534(.A1(new_n604), .A2(new_n233), .A3(new_n699), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n730), .B2(new_n512), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n729), .A2(KEYINPUT110), .A3(new_n575), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(G36gat), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n604), .A2(new_n735), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n512), .A2(G36gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n746), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n747), .A3(new_n750), .ZN(G1329gat));
  NAND3_X1  g550(.A1(new_n744), .A2(new_n241), .A3(new_n710), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n721), .A2(new_n558), .A3(new_n726), .A4(new_n728), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G43gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n754), .A3(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n757), .A3(G43gat), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n756), .A2(new_n758), .A3(new_n752), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(G1330gat));
  AOI21_X1  g560(.A(new_n242), .B1(new_n729), .B2(new_n356), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n743), .A2(G50gat), .A3(new_n355), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n762), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  INV_X1    g566(.A(new_n672), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n297), .A3(new_n642), .A4(new_n693), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n521), .A2(new_n551), .A3(new_n594), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n603), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n699), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n575), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT49), .B(G64gat), .Z(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1333gat));
  AND2_X1   g576(.A1(new_n771), .A2(new_n710), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n778), .A2(KEYINPUT113), .ZN(new_n779));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(KEYINPUT113), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n771), .A2(G71gat), .A3(new_n558), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g584(.A1(new_n771), .A2(new_n356), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT114), .B(G78gat), .Z(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n768), .A2(new_n296), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n693), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n721), .A2(new_n726), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n731), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n643), .B(new_n789), .C1(new_n723), .C2(new_n724), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n603), .A2(new_n770), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(KEYINPUT51), .A3(new_n643), .A4(new_n789), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n794), .A2(KEYINPUT115), .A3(new_n795), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n693), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n699), .A2(new_n613), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n793), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NAND4_X1  g603(.A1(new_n721), .A2(new_n575), .A3(new_n726), .A4(new_n791), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(G92gat), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n512), .A2(G92gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n733), .B(new_n808), .C1(new_n796), .C2(new_n799), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n614), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n802), .B2(new_n808), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n813), .B2(new_n815), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n792), .B2(new_n551), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n599), .A2(G99gat), .A3(new_n733), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT117), .Z(new_n819));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n721), .A2(new_n356), .A3(new_n726), .A4(new_n791), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n355), .A2(G106gat), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n800), .A2(new_n693), .A3(new_n801), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n796), .A2(new_n799), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n355), .A2(G106gat), .A3(new_n733), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT118), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n823), .A2(new_n826), .A3(new_n824), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n822), .A2(G106gat), .B1(new_n828), .B2(new_n829), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n824), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(G1339gat));
  NAND2_X1  g636(.A1(new_n694), .A2(new_n297), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n679), .A2(new_n680), .A3(new_n675), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n682), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n689), .B1(new_n681), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n692), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n848), .B(KEYINPUT55), .C1(new_n840), .C2(new_n842), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n286), .B(new_n213), .C1(new_n290), .C2(new_n292), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n206), .A2(new_n210), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n274), .A2(new_n275), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n262), .B1(new_n853), .B2(new_n261), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n285), .A2(new_n279), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n850), .A2(new_n642), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n851), .A2(new_n693), .A3(new_n856), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n297), .B2(new_n850), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n642), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n838), .B1(new_n861), .B2(new_n727), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n355), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n710), .A3(new_n699), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n575), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n296), .ZN(new_n866));
  MUX2_X1   g665(.A(new_n381), .B(G113gat), .S(new_n866), .Z(G1340gat));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n693), .ZN(new_n868));
  XNOR2_X1  g667(.A(KEYINPUT120), .B(G120gat), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1341gat));
  INV_X1    g669(.A(new_n865), .ZN(new_n871));
  INV_X1    g670(.A(new_n727), .ZN(new_n872));
  OAI21_X1  g671(.A(G127gat), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n865), .A2(new_n367), .A3(new_n768), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1342gat));
  NAND2_X1  g674(.A1(new_n643), .A2(new_n512), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT121), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n864), .A2(G134gat), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n864), .B2(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  NAND3_X1  g681(.A1(new_n699), .A2(new_n512), .A3(new_n551), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n679), .A2(new_n680), .A3(new_n675), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n681), .A3(new_n841), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n679), .A2(new_n680), .ZN(new_n886));
  INV_X1    g685(.A(new_n675), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n841), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n690), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n846), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n692), .A3(new_n843), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n296), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT122), .A3(new_n859), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n294), .B2(new_n295), .ZN(new_n896));
  INV_X1    g695(.A(new_n859), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n898), .A3(new_n642), .ZN(new_n899));
  INV_X1    g698(.A(new_n858), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n768), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n838), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT57), .B(new_n356), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n862), .A2(new_n356), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n903), .A2(KEYINPUT123), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n893), .A2(new_n859), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n643), .B1(new_n907), .B2(new_n895), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n858), .B1(new_n908), .B2(new_n894), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n838), .B1(new_n909), .B2(new_n768), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT57), .A4(new_n356), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n883), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n310), .B1(new_n913), .B2(new_n296), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n904), .A2(new_n883), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n310), .A3(new_n296), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n914), .A2(KEYINPUT58), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT58), .B1(new_n914), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1344gat));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n910), .B2(new_n356), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n356), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n693), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n924), .B2(new_n883), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n307), .A2(KEYINPUT59), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT124), .B(new_n928), .C1(new_n913), .C2(new_n693), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n906), .A2(new_n912), .ZN(new_n931));
  INV_X1    g730(.A(new_n883), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n693), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n926), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n307), .A3(new_n693), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1345gat));
  NAND3_X1  g736(.A1(new_n915), .A2(new_n314), .A3(new_n768), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n913), .A2(new_n727), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n314), .ZN(G1346gat));
  NAND2_X1  g739(.A1(new_n699), .A2(new_n551), .ZN(new_n941));
  OR4_X1    g740(.A1(G162gat), .A2(new_n904), .A3(new_n877), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n913), .A2(new_n643), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n315), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n699), .A2(new_n512), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n863), .A2(new_n710), .A3(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n946), .A2(new_n207), .A3(new_n297), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n945), .A2(new_n862), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(new_n596), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT125), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n296), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n951), .B2(new_n207), .ZN(G1348gat));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n457), .A3(new_n693), .ZN(new_n953));
  OAI21_X1  g752(.A(G176gat), .B1(new_n946), .B2(new_n733), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1349gat));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n464), .A3(new_n768), .ZN(new_n956));
  OAI21_X1  g755(.A(G183gat), .B1(new_n946), .B2(new_n872), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n956), .A2(new_n957), .B1(KEYINPUT126), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n959), .B(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n950), .A2(new_n465), .A3(new_n643), .ZN(new_n962));
  OAI21_X1  g761(.A(G190gat), .B1(new_n946), .B2(new_n642), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1351gat));
  NOR2_X1   g764(.A1(new_n558), .A2(new_n355), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n948), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n296), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n945), .A2(new_n551), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n899), .A2(new_n900), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n902), .B1(new_n971), .B2(new_n672), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n905), .B1(new_n972), .B2(new_n355), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n970), .B1(new_n973), .B2(new_n922), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n297), .A2(new_n209), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  NOR3_X1   g775(.A1(new_n967), .A2(G204gat), .A3(new_n733), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  OAI21_X1  g777(.A(G204gat), .B1(new_n924), .B2(new_n970), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1353gat));
  NAND3_X1  g779(.A1(new_n968), .A2(new_n300), .A3(new_n768), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  AOI211_X1 g781(.A(new_n982), .B(new_n300), .C1(new_n974), .C2(new_n768), .ZN(new_n983));
  INV_X1    g782(.A(new_n970), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n768), .B(new_n984), .C1(new_n921), .C2(new_n923), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g788(.A(KEYINPUT127), .B(new_n981), .C1(new_n983), .C2(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(G218gat), .B1(new_n968), .B2(new_n643), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n642), .A2(new_n301), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n974), .B2(new_n993), .ZN(G1355gat));
endmodule


