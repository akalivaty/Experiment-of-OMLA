//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(KEYINPUT64), .A3(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n195), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n198), .A2(KEYINPUT67), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(KEYINPUT67), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n192), .A2(new_n197), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT68), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(G128), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(G143), .B2(new_n191), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n205), .B(KEYINPUT68), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n200), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G104), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G107), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n214), .A3(G104), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(new_n217), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(KEYINPUT81), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n221), .A2(new_n222), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n220), .A3(new_n217), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n225), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT82), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n218), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT85), .B1(new_n212), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n218), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n227), .A2(new_n220), .A3(new_n217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n222), .B1(new_n235), .B2(new_n226), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n229), .A2(KEYINPUT82), .A3(new_n230), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n239));
  INV_X1    g053(.A(new_n200), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n243), .B2(new_n210), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n198), .B2(new_n209), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n200), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n232), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n233), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT66), .A2(G131), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G134), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n255), .B2(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(G134), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(new_n258), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n252), .B(new_n257), .C1(new_n260), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n263), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n254), .A2(new_n256), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n251), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n271), .A2(KEYINPUT86), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(KEYINPUT86), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n229), .A2(G101), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT4), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n228), .B2(new_n231), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT0), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n198), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n198), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n205), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n194), .A2(new_n279), .A3(new_n195), .A4(new_n197), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n229), .A2(new_n285), .A3(G101), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT83), .B1(new_n277), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT4), .B(new_n275), .C1(new_n236), .C2(new_n237), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT83), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n286), .A2(new_n283), .A3(new_n282), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n238), .A2(KEYINPUT84), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n232), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n296), .A4(new_n212), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n249), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n297), .A3(new_n268), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n250), .A2(KEYINPUT86), .A3(new_n271), .A4(new_n269), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n274), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT73), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G227), .ZN(new_n308));
  XOR2_X1   g122(.A(G110), .B(G140), .Z(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n288), .A2(new_n292), .B1(new_n298), .B2(new_n249), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n268), .B1(new_n313), .B2(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n302), .A2(new_n310), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G469), .B1(new_n316), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n300), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(new_n318), .B2(new_n314), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n274), .A2(new_n311), .A3(new_n300), .A4(new_n301), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G469), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n187), .B(new_n190), .C1(new_n317), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(G469), .A2(G902), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n302), .A2(new_n310), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n312), .A2(new_n315), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G469), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT87), .B1(new_n330), .B2(new_n189), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G475), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n340), .B2(new_n334), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(new_n191), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT72), .A2(G237), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT72), .A2(G237), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n307), .A2(new_n346), .A3(G143), .A4(G214), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n304), .B(new_n306), .C1(new_n344), .C2(new_n345), .ZN(new_n348));
  INV_X1    g162(.A(G214), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n196), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n342), .B1(KEYINPUT17), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n347), .A2(new_n350), .A3(new_n343), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n347), .A2(new_n350), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n358), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n347), .A2(new_n350), .A3(KEYINPUT91), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n340), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n191), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT79), .A4(new_n191), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n340), .A2(G146), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G113), .B(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(new_n216), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n357), .A2(new_n375), .A3(new_n378), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n333), .B1(new_n382), .B2(new_n323), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n357), .A2(new_n375), .A3(new_n378), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n353), .A2(new_n355), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n366), .A2(new_n367), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n340), .A2(KEYINPUT19), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n191), .A3(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n341), .A2(new_n191), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n364), .A2(new_n374), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n378), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n361), .A2(new_n363), .B1(new_n372), .B2(new_n373), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n391), .B1(new_n353), .B2(new_n355), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT92), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n384), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(G475), .A2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n385), .A2(new_n392), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n375), .A2(new_n403), .A3(new_n394), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n404), .A3(new_n379), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n381), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n400), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n383), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(G116), .ZN(new_n412));
  INV_X1    g226(.A(G116), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT93), .A3(G122), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(G116), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n214), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n207), .A2(G143), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n198), .A2(G143), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G134), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n255), .A3(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n415), .A2(KEYINPUT14), .B1(G116), .B2(new_n411), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(KEYINPUT14), .B2(new_n415), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G107), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n420), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n421), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n419), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G134), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n415), .A2(new_n416), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G107), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n417), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n424), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n419), .A2(KEYINPUT95), .A3(new_n255), .A4(new_n421), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n435), .A2(new_n438), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n429), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G217), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n188), .A2(new_n444), .A3(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n429), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n446), .A2(KEYINPUT96), .A3(new_n323), .A4(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G478), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(KEYINPUT15), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n409), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G119), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT2), .B(G113), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n289), .A2(new_n457), .A3(new_n286), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n294), .A2(new_n296), .ZN(new_n459));
  INV_X1    g273(.A(new_n454), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n413), .A2(KEYINPUT5), .A3(G119), .ZN(new_n463));
  INV_X1    g277(.A(G113), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n458), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n458), .C1(new_n459), .C2(new_n467), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n474), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n284), .A2(G125), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n244), .B2(G125), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n303), .A2(G224), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n469), .B(KEYINPUT8), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n238), .B2(new_n466), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n238), .B2(new_n466), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n477), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT7), .A3(new_n478), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n478), .A2(KEYINPUT7), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n477), .B(new_n488), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n490), .B2(new_n472), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT89), .Z(new_n494));
  XOR2_X1   g308(.A(new_n494), .B(KEYINPUT90), .Z(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n494), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n501), .A2(G952), .A3(new_n303), .ZN(new_n502));
  INV_X1    g316(.A(new_n307), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n503), .A2(G902), .A3(new_n501), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT21), .B(G898), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n499), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n332), .A2(new_n453), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n207), .A2(G119), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(G119), .B2(new_n198), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT24), .B(G110), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n514));
  INV_X1    g328(.A(G119), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(G128), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT77), .B(G110), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n390), .A3(new_n372), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(G110), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n342), .B(new_n522), .C1(new_n511), .C2(new_n512), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G137), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n523), .A3(new_n527), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G217), .A2(G902), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n444), .B2(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT75), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n323), .A3(new_n530), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(KEYINPUT25), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n534), .B(KEYINPUT76), .Z(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n537), .B2(KEYINPUT25), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT80), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT74), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n284), .B1(new_n264), .B2(new_n267), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n261), .A2(new_n256), .A3(G131), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n262), .B1(new_n261), .B2(new_n258), .ZN(new_n548));
  AOI211_X1 g362(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n253), .C2(G134), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n266), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n550), .B2(new_n343), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n545), .B(new_n456), .C1(new_n244), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n546), .B1(new_n557), .B2(G131), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n212), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n456), .A4(new_n545), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n244), .A2(new_n551), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n282), .A2(new_n283), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n550), .A2(new_n252), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n557), .A2(new_n251), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n457), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n555), .B1(new_n568), .B2(KEYINPUT28), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n307), .A2(new_n346), .A3(G210), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT27), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT29), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n556), .A2(new_n561), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT30), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n576), .A2(KEYINPUT69), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(KEYINPUT69), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n577), .B(new_n578), .C1(new_n562), .C2(new_n566), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n559), .A2(KEYINPUT69), .A3(new_n576), .A4(new_n545), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n457), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT70), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(new_n457), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n575), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n574), .B1(new_n586), .B2(new_n573), .ZN(new_n587));
  INV_X1    g401(.A(new_n573), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n588), .B(new_n555), .C1(new_n568), .C2(KEYINPUT28), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n589), .B2(KEYINPUT29), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n544), .B1(new_n591), .B2(G472), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT74), .B(new_n593), .C1(new_n587), .C2(new_n590), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n568), .A2(KEYINPUT28), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n554), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n588), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  INV_X1    g413(.A(new_n575), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n584), .B1(new_n581), .B2(new_n457), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT70), .B(new_n456), .C1(new_n579), .C2(new_n580), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n573), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n583), .A2(new_n585), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(KEYINPUT31), .A3(new_n573), .A4(new_n600), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n604), .A2(new_n593), .A3(new_n323), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT32), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n323), .B1(new_n603), .B2(new_n599), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT32), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n593), .A4(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n543), .B1(new_n595), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n509), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n230), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n618), .B2(new_n609), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n607), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n542), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n617), .B1(new_n622), .B2(new_n332), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n330), .A2(new_n189), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n187), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n330), .A2(KEYINPUT87), .A3(new_n189), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n627), .A2(KEYINPUT97), .A3(new_n542), .A4(new_n621), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n480), .A2(new_n491), .A3(new_n497), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n497), .B1(new_n480), .B2(new_n491), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n500), .B(new_n507), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n383), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n407), .B1(new_n406), .B2(new_n400), .ZN(new_n633));
  AOI211_X1 g447(.A(KEYINPUT20), .B(new_n401), .C1(new_n405), .C2(new_n381), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n446), .A2(new_n323), .A3(new_n448), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT100), .B1(new_n637), .B2(G478), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n639), .A3(new_n450), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n445), .A2(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n443), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT33), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n443), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT99), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n443), .B2(new_n642), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n648), .B(new_n649), .C1(new_n443), .C2(new_n642), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n446), .A2(new_n647), .A3(new_n448), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n450), .A2(G902), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n641), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n635), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n623), .A2(new_n628), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(new_n500), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n492), .A2(new_n494), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n498), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n635), .A2(new_n452), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT101), .A4(new_n507), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  INV_X1    g480(.A(new_n452), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n409), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n666), .B1(new_n631), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n623), .A2(new_n628), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n524), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n535), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n538), .B2(new_n540), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n620), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n509), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(new_n594), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n591), .A2(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT74), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n613), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n504), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n502), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n663), .A2(new_n664), .A3(new_n677), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n686), .A2(new_n627), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XNOR2_X1  g508(.A(new_n499), .B(KEYINPUT38), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n409), .A2(new_n452), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n500), .A3(new_n678), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n586), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n573), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n323), .B1(new_n568), .B2(new_n573), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n613), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n689), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n627), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT40), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n196), .ZN(G45));
  AND3_X1   g525(.A1(new_n646), .A2(new_n650), .A3(new_n651), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n712), .A2(new_n653), .B1(new_n638), .B2(new_n640), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n409), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n663), .A3(new_n677), .A4(new_n690), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n686), .A2(new_n627), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n321), .A2(new_n323), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n324), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(KEYINPUT103), .A3(G469), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n190), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n657), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n614), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n614), .A2(new_n670), .A3(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  OAI21_X1  g544(.A(new_n500), .B1(new_n629), .B2(new_n630), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n190), .B(new_n731), .C1(new_n722), .C2(new_n723), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n453), .A2(new_n506), .A3(new_n678), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n686), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  XNOR2_X1  g549(.A(new_n541), .B(KEYINPUT104), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n619), .A3(new_n607), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n696), .A2(new_n663), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n506), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n724), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR3_X1   g555(.A1(new_n409), .A2(new_n713), .A3(new_n689), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n679), .A2(new_n663), .A3(new_n742), .A4(new_n724), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  AND2_X1   g558(.A1(new_n686), .A2(new_n736), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n714), .A2(new_n690), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  INV_X1    g561(.A(new_n330), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n496), .A2(new_n189), .A3(new_n498), .A4(new_n500), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n495), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n480), .B2(new_n491), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n629), .A2(new_n752), .A3(new_n661), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT105), .A3(new_n189), .A4(new_n330), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n746), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n614), .A2(new_n755), .A3(KEYINPUT106), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT106), .B1(new_n614), .B2(new_n755), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND2_X1  g576(.A1(new_n750), .A2(new_n754), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n409), .A2(new_n667), .A3(new_n690), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n614), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  AND2_X1   g581(.A1(new_n316), .A2(KEYINPUT45), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n316), .B2(KEYINPUT45), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n326), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n326), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n324), .A3(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n189), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n777), .A3(new_n707), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n777), .B1(new_n776), .B2(new_n707), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n409), .A2(new_n655), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT43), .Z(new_n782));
  AND3_X1   g596(.A1(new_n782), .A2(new_n620), .A3(new_n677), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT44), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n753), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n780), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n253), .ZN(G39));
  XNOR2_X1  g601(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n776), .B(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n753), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n686), .A2(new_n542), .A3(new_n746), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT110), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(KEYINPUT111), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT112), .B(G140), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n722), .A2(new_n723), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n190), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n782), .A2(new_n502), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n621), .A3(new_n736), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(new_n791), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n695), .A2(new_n500), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n724), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n724), .A2(new_n753), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT117), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n542), .A2(new_n813), .A3(new_n502), .A4(new_n704), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n409), .A3(new_n713), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n813), .A2(new_n804), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n679), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n801), .B1(new_n807), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n732), .ZN(new_n820));
  OAI211_X1 g634(.A(G952), .B(new_n303), .C1(new_n805), .C2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n814), .B2(new_n714), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n745), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT48), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n816), .A2(KEYINPUT48), .A3(new_n745), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n818), .B(KEYINPUT118), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT51), .B1(new_n803), .B2(new_n806), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n819), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n689), .A2(new_n190), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n676), .B(new_n832), .C1(new_n538), .C2(new_n540), .ZN(new_n833));
  AOI211_X1 g647(.A(KEYINPUT114), .B(new_n833), .C1(new_n317), .C2(new_n324), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n835));
  INV_X1    g649(.A(new_n833), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n330), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n738), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n703), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n693), .A2(new_n717), .A3(new_n840), .A4(new_n743), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n715), .B1(new_n595), .B2(new_n613), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n738), .B1(new_n613), .B2(new_n702), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n844), .A2(new_n627), .B1(new_n845), .B2(new_n838), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n691), .B1(new_n595), .B2(new_n613), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n607), .A2(new_n742), .A3(new_n619), .A4(new_n677), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n627), .B1(new_n848), .B2(new_n732), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n842), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n843), .B1(new_n842), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n729), .A2(new_n726), .A3(new_n734), .A4(new_n740), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n791), .A2(new_n453), .A3(new_n678), .A4(new_n689), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n686), .A3(new_n627), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n763), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n766), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n664), .A2(KEYINPUT113), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT113), .B1(new_n714), .B2(new_n664), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n508), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n623), .A2(new_n628), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n509), .B1(new_n614), .B2(new_n679), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n860), .A2(new_n761), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n831), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n614), .A2(new_n725), .B1(new_n739), .B2(new_n724), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n729), .A4(new_n734), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n761), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n859), .A2(new_n831), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n866), .A2(new_n876), .A3(new_n851), .A4(new_n842), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n869), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT53), .B1(new_n854), .B2(new_n867), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n860), .A2(new_n761), .A3(new_n866), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n831), .A3(new_n851), .A4(new_n842), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n879), .B1(new_n883), .B2(new_n869), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n830), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n736), .A2(new_n189), .A3(new_n500), .ZN(new_n886));
  OR4_X1    g700(.A1(new_n703), .A2(new_n695), .A3(new_n781), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n802), .B(KEYINPUT49), .Z(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n307), .A2(G952), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n473), .A2(new_n475), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n479), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n878), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(G902), .A3(new_n494), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(G902), .A3(new_n495), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n897), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n900), .B2(new_n894), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n890), .B(new_n898), .C1(new_n899), .C2(new_n902), .ZN(G51));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n770), .B(KEYINPUT121), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n841), .A2(KEYINPUT52), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n850), .B1(new_n846), .B2(new_n849), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT115), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n842), .A2(new_n851), .A3(new_n843), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT53), .B1(new_n910), .B2(new_n881), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n875), .A2(new_n877), .ZN(new_n912));
  OAI211_X1 g726(.A(G902), .B(new_n905), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n326), .B(KEYINPUT57), .Z(new_n915));
  AOI21_X1  g729(.A(new_n869), .B1(new_n868), .B2(new_n878), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n911), .A2(KEYINPUT54), .A3(new_n912), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n918), .B2(new_n321), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n904), .B1(new_n919), .B2(new_n890), .ZN(new_n920));
  INV_X1    g734(.A(new_n890), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n879), .A2(new_n922), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n923), .A2(new_n915), .B1(new_n319), .B2(new_n320), .ZN(new_n924));
  OAI211_X1 g738(.A(KEYINPUT122), .B(new_n921), .C1(new_n924), .C2(new_n914), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G54));
  NAND2_X1  g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n895), .A2(G902), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n399), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n895), .A2(G902), .A3(new_n406), .A4(new_n928), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n921), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n921), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G60));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT59), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n923), .A2(new_n712), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n712), .B1(new_n884), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n890), .ZN(G63));
  XNOR2_X1  g755(.A(new_n532), .B(KEYINPUT60), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n868), .B2(new_n878), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n531), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n890), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n675), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n945), .A2(KEYINPUT124), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n947), .B(new_n921), .C1(new_n531), .C2(new_n943), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n948), .A2(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n505), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n866), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n855), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n957), .B2(new_n503), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n891), .B1(G898), .B2(new_n307), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n958), .B(new_n960), .ZN(G69));
  AOI21_X1  g775(.A(new_n786), .B1(new_n796), .B2(new_n797), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n839), .B(new_n745), .C1(new_n778), .C2(new_n779), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n849), .A2(new_n717), .A3(new_n766), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n963), .A2(new_n761), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n965), .A3(new_n307), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n387), .A2(new_n388), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n581), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n503), .A2(G900), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n791), .B1(new_n861), .B2(new_n862), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n614), .A2(new_n971), .A3(new_n627), .A4(new_n707), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n849), .A2(new_n717), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n710), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n503), .B1(new_n978), .B2(new_n962), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(new_n968), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n307), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n970), .B(new_n983), .C1(new_n979), .C2(new_n968), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(new_n586), .A2(new_n588), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT127), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n962), .A2(new_n957), .A3(new_n965), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n699), .A2(new_n990), .A3(new_n986), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n883), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n994), .A3(new_n921), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n978), .A2(new_n957), .A3(new_n962), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n699), .B1(new_n996), .B2(new_n990), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(G57));
endmodule


