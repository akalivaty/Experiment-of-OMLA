//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT69), .A3(G116), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n192), .C1(G116), .C2(new_n191), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT30), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT68), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(KEYINPUT68), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT67), .B1(new_n210), .B2(new_n205), .ZN(new_n211));
  AND4_X1   g025(.A1(KEYINPUT67), .A2(new_n205), .A3(new_n201), .A4(new_n207), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n203), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT11), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n219), .A2(KEYINPUT11), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n219), .A2(KEYINPUT11), .A3(G134), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n222), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n219), .B2(G134), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n214), .A2(KEYINPUT66), .A3(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n201), .A2(new_n207), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT0), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n204), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n210), .A2(KEYINPUT0), .A3(G128), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n223), .B1(new_n218), .B2(new_n220), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n222), .B1(new_n244), .B2(new_n226), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n215), .A2(new_n217), .B1(KEYINPUT11), .B2(new_n219), .ZN(new_n246));
  NOR4_X1   g060(.A1(new_n246), .A2(G131), .A3(new_n225), .A4(new_n223), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n197), .B(new_n199), .C1(new_n234), .C2(new_n248), .ZN(new_n249));
  AND4_X1   g063(.A1(KEYINPUT68), .A2(new_n234), .A3(new_n248), .A4(new_n196), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n195), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT31), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(G101), .ZN(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n254), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n234), .A2(new_n248), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n195), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n251), .A2(new_n252), .A3(new_n258), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g077(.A(new_n258), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(new_n195), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n234), .A2(new_n248), .A3(KEYINPUT72), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT72), .B1(new_n234), .B2(new_n248), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n259), .A2(new_n195), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n261), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n264), .B(new_n269), .C1(new_n271), .C2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(new_n197), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n205), .A2(new_n201), .A3(new_n207), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n210), .A2(KEYINPUT67), .A3(new_n205), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n202), .B(new_n208), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n227), .A2(new_n233), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n241), .A2(new_n242), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n221), .A2(new_n224), .A3(new_n226), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G131), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n227), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n273), .B(new_n198), .C1(new_n280), .C2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n234), .A2(new_n248), .A3(KEYINPUT68), .A4(new_n196), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n260), .B1(new_n287), .B2(new_n195), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n252), .A4(new_n258), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n263), .A2(new_n272), .A3(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n264), .B(new_n260), .C1(new_n287), .C2(new_n195), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT70), .B1(new_n292), .B2(new_n252), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n251), .A2(new_n258), .A3(new_n261), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT31), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT73), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  INV_X1    g115(.A(new_n299), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n301), .B(new_n302), .C1(new_n291), .C2(new_n297), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n291), .B2(new_n297), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n269), .B1(new_n271), .B2(new_n265), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n306), .B2(new_n258), .ZN(new_n307));
  INV_X1    g121(.A(new_n288), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n264), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(KEYINPUT29), .A3(new_n258), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n305), .A2(KEYINPUT32), .B1(new_n313), .B2(G472), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(G110), .B(G122), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT87), .B(KEYINPUT8), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  INV_X1    g134(.A(G104), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(G107), .ZN(new_n322));
  INV_X1    g136(.A(G107), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT3), .A3(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(G107), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT79), .B(G101), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n319), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n322), .A2(new_n324), .B1(new_n321), .B2(G107), .ZN(new_n330));
  INV_X1    g144(.A(new_n328), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(KEYINPUT80), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(KEYINPUT82), .A3(G107), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(new_n335), .C1(new_n321), .C2(G107), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n329), .A2(new_n332), .B1(G101), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n191), .A3(G116), .ZN(new_n339));
  OAI211_X1 g153(.A(G113), .B(new_n339), .C1(new_n193), .C2(new_n338), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n193), .A2(new_n194), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n337), .A2(new_n342), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n318), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n327), .A2(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(new_n332), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n327), .A2(KEYINPUT81), .A3(KEYINPUT4), .A4(G101), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n195), .ZN(new_n354));
  INV_X1    g168(.A(new_n316), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n343), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT86), .B1(new_n243), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n281), .A2(new_n359), .A3(G125), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G224), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(G953), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n278), .A2(new_n357), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(KEYINPUT7), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n358), .A3(new_n360), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT7), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n346), .A2(new_n356), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n311), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n316), .B(KEYINPUT85), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n354), .B2(new_n343), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT6), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n354), .A2(new_n343), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n356), .B1(new_n376), .B2(new_n373), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(KEYINPUT6), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n367), .B(new_n364), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G210), .B1(G237), .B2(G902), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n372), .B(new_n381), .C1(new_n378), .C2(new_n379), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n256), .A2(G952), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(G234), .B2(G237), .ZN(new_n390));
  INV_X1    g204(.A(G234), .ZN(new_n391));
  OAI211_X1 g205(.A(G902), .B(G953), .C1(new_n391), .C2(new_n255), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n392), .B(KEYINPUT92), .Z(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT21), .B(G898), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n200), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n255), .A2(new_n256), .A3(G214), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n206), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(G131), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n401), .B(G143), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n222), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n400), .B(new_n403), .C1(new_n407), .C2(KEYINPUT17), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n321), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n405), .B1(new_n411), .B2(new_n222), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n398), .B(new_n200), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n412), .B(new_n413), .C1(new_n411), .C2(new_n404), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n398), .B2(KEYINPUT89), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n398), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT19), .B1(new_n420), .B2(KEYINPUT88), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n421), .B2(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n200), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n399), .A2(G146), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n407), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n425), .A2(new_n414), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n415), .B1(new_n426), .B2(new_n410), .ZN(new_n427));
  INV_X1    g241(.A(G475), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n427), .A2(KEYINPUT20), .A3(new_n428), .A4(new_n311), .ZN(new_n429));
  INV_X1    g243(.A(new_n415), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n410), .B1(new_n425), .B2(new_n414), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n428), .B(new_n311), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n410), .B1(new_n408), .B2(new_n414), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n311), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G475), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n218), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G122), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(new_n323), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n323), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n446));
  OR3_X1    g260(.A1(new_n204), .A2(KEYINPUT13), .A3(G143), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n446), .A2(G134), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT90), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n442), .B(new_n323), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(G134), .A3(new_n447), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n441), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n218), .A2(new_n440), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n323), .B1(new_n459), .B2(KEYINPUT14), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n455), .A2(new_n441), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n443), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT9), .B(G234), .Z(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(G217), .A3(new_n256), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n454), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n454), .B2(new_n463), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n311), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(KEYINPUT15), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(KEYINPUT91), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n311), .C1(new_n467), .C2(new_n468), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AND4_X1   g291(.A1(new_n396), .A2(new_n439), .A3(new_n472), .A4(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n388), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(KEYINPUT24), .B(G110), .Z(new_n480));
  NAND2_X1  g294(.A1(new_n191), .A2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n204), .A2(G119), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n400), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G110), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(KEYINPUT23), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n204), .A3(G119), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(new_n481), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT75), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n489), .A2(new_n485), .A3(new_n481), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n494));
  OAI221_X1 g308(.A(new_n424), .B1(G146), .B2(new_n420), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(G137), .ZN(new_n498));
  INV_X1    g312(.A(G221), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n499), .A2(new_n391), .A3(G953), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n498), .B(new_n500), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n492), .A2(new_n495), .A3(new_n501), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G217), .B1(new_n391), .B2(G902), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT74), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n311), .ZN(new_n508));
  XOR2_X1   g322(.A(new_n508), .B(KEYINPUT78), .Z(new_n509));
  NOR2_X1   g323(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n511));
  OR3_X1    g325(.A1(new_n505), .A2(G902), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n505), .B2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n499), .B1(new_n464), .B2(new_n311), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G140), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n256), .A2(G227), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  NAND2_X1  g336(.A1(new_n353), .A2(new_n243), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n336), .A2(G101), .ZN(new_n526));
  INV_X1    g340(.A(new_n332), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT80), .B1(new_n330), .B2(new_n331), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n529), .B2(new_n278), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n245), .A2(new_n247), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(KEYINPUT84), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n523), .A2(new_n532), .A3(new_n530), .A4(new_n524), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n529), .A2(new_n278), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n337), .A2(new_n213), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n533), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n337), .B(new_n213), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(new_n544), .A3(new_n545), .A4(new_n533), .ZN(new_n550));
  AND4_X1   g364(.A1(new_n539), .A2(new_n548), .A3(new_n522), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n519), .B(new_n311), .C1(new_n540), .C2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n539), .A2(new_n522), .ZN(new_n553));
  INV_X1    g367(.A(new_n522), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n550), .A3(new_n539), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n538), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G469), .B1(new_n556), .B2(G902), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n518), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n315), .A2(new_n479), .A3(new_n517), .A4(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n328), .ZN(G3));
  AOI211_X1 g374(.A(KEYINPUT70), .B(new_n252), .C1(new_n288), .C2(new_n258), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n295), .B1(new_n294), .B2(KEYINPUT31), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n263), .A2(new_n272), .A3(new_n290), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n299), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n301), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n298), .A2(new_n311), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G472), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n517), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n552), .A2(new_n557), .ZN(new_n573));
  INV_X1    g387(.A(new_n518), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n384), .A2(KEYINPUT93), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n387), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n383), .A2(KEYINPUT93), .A3(new_n384), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n467), .B2(new_n468), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n454), .A2(new_n463), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT95), .B1(new_n583), .B2(new_n466), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(KEYINPUT33), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n467), .B2(new_n468), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n471), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n473), .A2(new_n471), .A3(new_n476), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n439), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n580), .A2(new_n395), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n576), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  AOI21_X1  g412(.A(new_n438), .B1(new_n477), .B2(new_n472), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n580), .A2(new_n395), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n576), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G107), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NAND2_X1  g418(.A1(new_n515), .A2(new_n516), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n496), .ZN(new_n607));
  INV_X1    g421(.A(new_n509), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n573), .A2(new_n574), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n479), .A2(new_n568), .A3(new_n570), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT37), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n485), .ZN(G12));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n578), .A2(new_n579), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT32), .B1(new_n566), .B2(new_n567), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n313), .A2(G472), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n611), .B(new_n616), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(G900), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n393), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n390), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n599), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n615), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n558), .A2(new_n610), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n304), .B2(new_n314), .ZN(new_n629));
  INV_X1    g443(.A(new_n626), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n616), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XNOR2_X1  g447(.A(new_n385), .B(KEYINPUT97), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT38), .ZN(new_n635));
  INV_X1    g449(.A(new_n618), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n288), .A2(new_n264), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n271), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n640), .B2(new_n264), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n617), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n643), .A2(new_n387), .A3(new_n610), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n439), .B1(new_n472), .B2(new_n477), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n625), .B(KEYINPUT39), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n558), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT40), .Z(new_n648));
  NAND4_X1  g462(.A1(new_n635), .A2(new_n644), .A3(new_n645), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  AND3_X1   g464(.A1(new_n591), .A2(new_n438), .A3(new_n625), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n578), .A2(new_n579), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n629), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  INV_X1    g470(.A(new_n537), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT84), .B1(new_n531), .B2(new_n533), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n539), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n551), .B1(new_n659), .B2(new_n554), .ZN(new_n660));
  OAI21_X1  g474(.A(G469), .B1(new_n660), .B2(G902), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n552), .A3(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(G469), .C1(new_n660), .C2(G902), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n574), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n315), .A3(new_n595), .A4(new_n517), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n315), .A3(new_n601), .A4(new_n517), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  INV_X1    g486(.A(new_n610), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n674), .A2(new_n478), .A3(new_n315), .A4(new_n616), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G119), .ZN(G21));
  NOR2_X1   g490(.A1(new_n666), .A2(new_n395), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n578), .A2(new_n579), .A3(new_n645), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n578), .A2(KEYINPUT101), .A3(new_n579), .A4(new_n645), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n569), .A2(new_n683), .A3(G472), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n292), .A2(new_n252), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n299), .B1(new_n564), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n291), .B2(new_n297), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT100), .B1(new_n687), .B2(new_n637), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n677), .A2(new_n682), .A3(new_n517), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT102), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n458), .ZN(G24));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n652), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G125), .ZN(G27));
  NOR2_X1   g510(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n517), .B1(new_n620), .B2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n651), .A2(new_n386), .A3(new_n383), .A4(new_n384), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n575), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n700), .B(new_n517), .C1(new_n617), .C2(new_n620), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n315), .A2(KEYINPUT103), .A3(new_n517), .A4(new_n700), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n702), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT104), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n706), .A2(new_n707), .A3(new_n710), .A4(new_n702), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n703), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n222), .ZN(G33));
  NOR2_X1   g527(.A1(new_n617), .A2(new_n620), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n572), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n383), .A2(new_n386), .A3(new_n384), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n715), .A2(new_n558), .A3(new_n630), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n214), .ZN(G36));
  AOI21_X1  g533(.A(new_n673), .B1(new_n568), .B2(new_n570), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n439), .A2(new_n591), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT43), .Z(new_n723));
  AND2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n556), .B(KEYINPUT45), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND2_X1  g542(.A1(G469), .A2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(G469), .C1(new_n727), .C2(G902), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n552), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n574), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n646), .B(new_n735), .C1(new_n724), .C2(KEYINPUT44), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT106), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G137), .ZN(G39));
  NOR2_X1   g553(.A1(new_n699), .A2(new_n517), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n734), .A2(new_n741), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n714), .B(new_n740), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G140), .ZN(G42));
  XOR2_X1   g560(.A(new_n665), .B(KEYINPUT49), .Z(new_n747));
  NAND2_X1  g561(.A1(new_n643), .A2(new_n517), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n439), .A2(new_n386), .A3(new_n591), .A4(new_n574), .ZN(new_n749));
  OR4_X1    g563(.A1(new_n635), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n667), .A2(new_n390), .A3(new_n717), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT111), .Z(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n439), .A3(new_n592), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n689), .A2(new_n624), .A3(new_n572), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n723), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n666), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n635), .A2(new_n386), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT50), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT50), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n744), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n665), .A2(new_n518), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n742), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n717), .A3(new_n723), .A4(new_n755), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n667), .A2(new_n723), .A3(new_n390), .A4(new_n717), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n766), .A2(new_n673), .A3(new_n689), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n754), .A2(new_n761), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n761), .A2(new_n770), .A3(new_n765), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n389), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n753), .A2(new_n593), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n766), .A2(new_n698), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT48), .Z(new_n778));
  NAND2_X1  g592(.A1(new_n757), .A2(new_n616), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n709), .A2(new_n711), .ZN(new_n783));
  INV_X1    g597(.A(new_n703), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n691), .A2(new_n675), .A3(new_n668), .A4(new_n671), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n654), .A2(new_n629), .B1(new_n674), .B2(new_n694), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n642), .B1(new_n568), .B2(new_n187), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n610), .B1(new_n788), .B2(new_n618), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n558), .A3(new_n625), .A4(new_n682), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n632), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n786), .B1(new_n791), .B2(KEYINPUT52), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n632), .A2(new_n787), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n785), .A2(new_n792), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n594), .A2(new_n600), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n576), .A2(new_n396), .A3(new_n388), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n559), .A3(new_n612), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n439), .A2(new_n472), .A3(new_n477), .A4(new_n625), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n716), .B2(new_n801), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n716), .A2(new_n801), .A3(new_n800), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n315), .A2(new_n558), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n690), .A2(new_n700), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n673), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n799), .A2(new_n718), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n785), .A2(new_n792), .A3(new_n795), .A4(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n796), .A2(new_n808), .A3(KEYINPUT53), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(KEYINPUT53), .B2(new_n796), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n781), .B(new_n782), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n795), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n712), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n792), .A4(new_n807), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT109), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n785), .A2(new_n792), .A3(new_n795), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n807), .C1(new_n793), .C2(new_n812), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n796), .A2(new_n808), .A3(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT54), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n811), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT110), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n811), .C1(new_n819), .C2(new_n823), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n780), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(G952), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n256), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT113), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n750), .B1(new_n828), .B2(new_n831), .ZN(G75));
  NAND4_X1  g646(.A1(new_n821), .A2(G210), .A3(G902), .A4(new_n822), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT114), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(G953), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT115), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n834), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n378), .B(new_n379), .Z(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT55), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n835), .B(new_n838), .C1(new_n842), .C2(new_n843), .ZN(G51));
  XNOR2_X1  g658(.A(new_n729), .B(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n782), .B1(new_n809), .B2(new_n810), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(KEYINPUT116), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n850), .A2(new_n851), .B1(new_n540), .B2(new_n551), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n728), .B(KEYINPUT117), .Z(new_n853));
  NAND4_X1  g667(.A1(new_n821), .A2(G902), .A3(new_n822), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n838), .B1(new_n852), .B2(new_n854), .ZN(G54));
  NAND4_X1  g669(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT58), .A4(G902), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n428), .ZN(new_n857));
  INV_X1    g671(.A(new_n427), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n856), .A2(new_n428), .A3(new_n427), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n837), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(KEYINPUT118), .B(new_n837), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(G60));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n866));
  NAND2_X1  g680(.A1(G478), .A2(G902), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n847), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n823), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n585), .A2(new_n587), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n837), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n825), .A2(new_n827), .A3(new_n868), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n871), .ZN(G63));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT121), .Z(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT60), .Z(new_n877));
  NAND4_X1  g691(.A1(new_n821), .A2(new_n822), .A3(new_n607), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n821), .A2(new_n822), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n505), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT123), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n882), .B2(KEYINPUT123), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n883), .A3(new_n837), .A4(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n880), .A2(new_n837), .A3(new_n882), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G66));
  NOR2_X1   g703(.A1(new_n786), .A2(new_n799), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(G953), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  OAI21_X1  g706(.A(G953), .B1(new_n394), .B2(new_n362), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n378), .B1(G898), .B2(new_n256), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(G69));
  NOR2_X1   g710(.A1(new_n256), .A2(G227), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n745), .B1(new_n726), .B2(new_n736), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n899));
  INV_X1    g713(.A(new_n647), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n715), .A2(new_n900), .A3(new_n717), .A4(new_n797), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n632), .A2(new_n787), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n649), .ZN(new_n903));
  NOR2_X1   g717(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n897), .B1(new_n906), .B2(new_n256), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n287), .B(new_n422), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n622), .B2(G953), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n897), .A2(G900), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n898), .A2(new_n718), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n698), .B1(new_n680), .B2(new_n681), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n735), .A2(new_n646), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n712), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n916), .B2(G953), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n907), .A2(new_n909), .B1(new_n917), .B2(new_n908), .ZN(G72));
  NAND2_X1  g732(.A1(G472), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT63), .Z(new_n920));
  NOR2_X1   g734(.A1(new_n308), .A2(new_n258), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n639), .A2(new_n817), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n899), .A2(new_n890), .A3(new_n901), .A4(new_n905), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n639), .B1(new_n924), .B2(new_n920), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n921), .B(KEYINPUT126), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n911), .A2(new_n890), .A3(new_n915), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n920), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n928), .A2(new_n929), .A3(new_n838), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n928), .B2(new_n838), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n923), .B(new_n925), .C1(new_n930), .C2(new_n931), .ZN(G57));
endmodule


