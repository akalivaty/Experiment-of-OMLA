

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U545 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X2 U546 ( .A1(G8), .A2(n711), .ZN(n761) );
  NAND2_X2 U547 ( .A1(n675), .A2(n674), .ZN(n711) );
  INV_X2 U548 ( .A(n711), .ZN(n706) );
  OR2_X1 U549 ( .A1(n721), .A2(n720), .ZN(n734) );
  BUF_X1 U550 ( .A(n672), .Z(G160) );
  XOR2_X1 U551 ( .A(KEYINPUT17), .B(n536), .Z(n884) );
  XNOR2_X1 U552 ( .A(n730), .B(KEYINPUT32), .ZN(n731) );
  XNOR2_X1 U553 ( .A(n732), .B(n731), .ZN(n753) );
  NOR2_X1 U554 ( .A1(G651), .A2(n619), .ZN(n627) );
  NOR2_X1 U555 ( .A1(G651), .A2(G543), .ZN(n632) );
  XOR2_X1 U556 ( .A(KEYINPUT0), .B(G543), .Z(n619) );
  NAND2_X1 U557 ( .A1(n627), .A2(G52), .ZN(n515) );
  XOR2_X1 U558 ( .A(G651), .B(KEYINPUT66), .Z(n517) );
  NOR2_X1 U559 ( .A1(G543), .A2(n517), .ZN(n513) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n513), .Z(n628) );
  NAND2_X1 U561 ( .A1(G64), .A2(n628), .ZN(n514) );
  NAND2_X1 U562 ( .A1(n515), .A2(n514), .ZN(n522) );
  NAND2_X1 U563 ( .A1(n632), .A2(G90), .ZN(n516) );
  XOR2_X1 U564 ( .A(KEYINPUT67), .B(n516), .Z(n519) );
  NOR2_X1 U565 ( .A1(n619), .A2(n517), .ZN(n633) );
  NAND2_X1 U566 ( .A1(G77), .A2(n633), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U568 ( .A(KEYINPUT9), .B(n520), .Z(n521) );
  NOR2_X1 U569 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT68), .B(n523), .Z(G301) );
  INV_X1 U571 ( .A(G301), .ZN(G171) );
  NAND2_X1 U572 ( .A1(n632), .A2(G91), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G78), .A2(n633), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U575 ( .A1(n627), .A2(G53), .ZN(n527) );
  NAND2_X1 U576 ( .A1(G65), .A2(n628), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n528) );
  OR2_X1 U578 ( .A1(n529), .A2(n528), .ZN(G299) );
  NAND2_X1 U579 ( .A1(n632), .A2(G85), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G72), .A2(n633), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n627), .A2(G47), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G60), .A2(n628), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n534) );
  OR2_X1 U585 ( .A1(n535), .A2(n534), .ZN(G290) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G137), .A2(n884), .ZN(n538) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U590 ( .A1(G113), .A2(n889), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U592 ( .A(n539), .B(KEYINPUT65), .ZN(n547) );
  INV_X1 U593 ( .A(G2104), .ZN(n540) );
  AND2_X1 U594 ( .A1(n540), .A2(G2105), .ZN(n891) );
  AND2_X1 U595 ( .A1(G125), .A2(n891), .ZN(n545) );
  INV_X1 U596 ( .A(KEYINPUT23), .ZN(n543) );
  NOR2_X1 U597 ( .A1(n540), .A2(G2105), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT64), .ZN(n885) );
  AND2_X1 U599 ( .A1(G101), .A2(n885), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n543), .B(n542), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  AND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n672) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  NAND2_X1 U606 ( .A1(n632), .A2(G89), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G76), .A2(n633), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT5), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n627), .A2(G51), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G63), .A2(n628), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n555), .Z(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U616 ( .A(n558), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U620 ( .A(G223), .B(KEYINPUT69), .ZN(n817) );
  NAND2_X1 U621 ( .A1(n817), .A2(G567), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U623 ( .A(G860), .B(KEYINPUT72), .Z(n584) );
  NAND2_X1 U624 ( .A1(G81), .A2(n632), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT70), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G68), .A2(n633), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(n565), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n628), .A2(G56), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n566), .Z(n569) );
  NAND2_X1 U632 ( .A1(G43), .A2(n627), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(n567), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n945) );
  OR2_X1 U636 ( .A1(n584), .A2(n945), .ZN(G153) );
  INV_X1 U637 ( .A(G868), .ZN(n647) );
  NOR2_X1 U638 ( .A1(n647), .A2(G171), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT73), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n627), .A2(G54), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G66), .A2(n628), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n632), .A2(G92), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G79), .A2(n633), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT15), .ZN(n940) );
  NAND2_X1 U648 ( .A1(n647), .A2(n940), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G284) );
  NOR2_X1 U650 ( .A1(G868), .A2(G299), .ZN(n583) );
  NOR2_X1 U651 ( .A1(G286), .A2(n647), .ZN(n582) );
  NOR2_X1 U652 ( .A1(n583), .A2(n582), .ZN(G297) );
  NAND2_X1 U653 ( .A1(n584), .A2(G559), .ZN(n585) );
  INV_X1 U654 ( .A(n940), .ZN(n901) );
  NAND2_X1 U655 ( .A1(n585), .A2(n901), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U657 ( .A1(G868), .A2(n945), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G868), .A2(n901), .ZN(n587) );
  NOR2_X1 U659 ( .A1(G559), .A2(n587), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(G282) );
  NAND2_X1 U661 ( .A1(G111), .A2(n889), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT74), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n885), .A2(G99), .ZN(n591) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n591), .Z(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G123), .A2(n891), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT18), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n884), .A2(G135), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n967) );
  XOR2_X1 U671 ( .A(G2096), .B(n967), .Z(n599) );
  NOR2_X1 U672 ( .A1(G2100), .A2(n599), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT76), .B(n600), .Z(G156) );
  NAND2_X1 U674 ( .A1(n628), .A2(G67), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT78), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G93), .A2(n632), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G55), .A2(n627), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G80), .A2(n633), .ZN(n604) );
  XNOR2_X1 U680 ( .A(KEYINPUT77), .B(n604), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n648) );
  NAND2_X1 U683 ( .A1(n901), .A2(G559), .ZN(n644) );
  XNOR2_X1 U684 ( .A(n945), .B(n644), .ZN(n609) );
  NOR2_X1 U685 ( .A1(G860), .A2(n609), .ZN(n610) );
  XOR2_X1 U686 ( .A(n648), .B(n610), .Z(G145) );
  NAND2_X1 U687 ( .A1(G86), .A2(n632), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G48), .A2(n627), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n633), .A2(G73), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT81), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT2), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G61), .A2(n628), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G305) );
  NAND2_X1 U696 ( .A1(G49), .A2(n627), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G87), .A2(n619), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n628), .A2(n622), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n623), .Z(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U703 ( .A(KEYINPUT80), .B(n626), .ZN(G288) );
  NAND2_X1 U704 ( .A1(n627), .A2(G50), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G62), .A2(n628), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT82), .B(n631), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n632), .A2(G88), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G75), .A2(n633), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(G166) );
  INV_X1 U712 ( .A(G166), .ZN(G303) );
  XOR2_X1 U713 ( .A(G290), .B(G299), .Z(n638) );
  XNOR2_X1 U714 ( .A(n648), .B(n638), .ZN(n639) );
  XNOR2_X1 U715 ( .A(KEYINPUT19), .B(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(G305), .B(G288), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n642), .B(G303), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n643), .B(n945), .ZN(n900) );
  XNOR2_X1 U720 ( .A(n900), .B(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n645), .A2(G868), .ZN(n646) );
  XOR2_X1 U722 ( .A(KEYINPUT83), .B(n646), .Z(n650) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(G295) );
  NAND2_X1 U725 ( .A1(G2084), .A2(G2078), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT20), .B(n651), .Z(n652) );
  NAND2_X1 U727 ( .A1(G2090), .A2(n652), .ZN(n653) );
  XNOR2_X1 U728 ( .A(KEYINPUT21), .B(n653), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n654), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U730 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U731 ( .A1(G220), .A2(G219), .ZN(n655) );
  XOR2_X1 U732 ( .A(KEYINPUT22), .B(n655), .Z(n656) );
  NOR2_X1 U733 ( .A1(G218), .A2(n656), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G96), .A2(n657), .ZN(n822) );
  NAND2_X1 U735 ( .A1(G2106), .A2(n822), .ZN(n661) );
  NAND2_X1 U736 ( .A1(G69), .A2(G120), .ZN(n658) );
  NOR2_X1 U737 ( .A1(G237), .A2(n658), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G108), .A2(n659), .ZN(n823) );
  NAND2_X1 U739 ( .A1(G567), .A2(n823), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n852) );
  NAND2_X1 U741 ( .A1(G661), .A2(G483), .ZN(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT84), .B(n662), .ZN(n663) );
  NOR2_X1 U743 ( .A1(n852), .A2(n663), .ZN(n821) );
  NAND2_X1 U744 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U745 ( .A1(G126), .A2(n891), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G114), .A2(n889), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n671) );
  INV_X1 U748 ( .A(KEYINPUT85), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n884), .A2(G138), .ZN(n667) );
  NAND2_X1 U750 ( .A1(G102), .A2(n885), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G164) );
  XNOR2_X1 U754 ( .A(G1986), .B(G290), .ZN(n950) );
  NAND2_X1 U755 ( .A1(n672), .A2(G40), .ZN(n673) );
  NOR2_X1 U756 ( .A1(G164), .A2(G1384), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n673), .A2(n674), .ZN(n812) );
  NAND2_X1 U758 ( .A1(n950), .A2(n812), .ZN(n801) );
  XNOR2_X1 U759 ( .A(n673), .B(KEYINPUT91), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n706), .A2(G2072), .ZN(n677) );
  INV_X1 U761 ( .A(KEYINPUT27), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n677), .B(n676), .ZN(n679) );
  INV_X1 U763 ( .A(n706), .ZN(n722) );
  NAND2_X1 U764 ( .A1(G1956), .A2(n722), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n700) );
  NOR2_X1 U766 ( .A1(G299), .A2(n700), .ZN(n680) );
  XNOR2_X1 U767 ( .A(n680), .B(KEYINPUT94), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G1348), .A2(n722), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G2067), .A2(n706), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U771 ( .A1(n940), .A2(n683), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n699) );
  NAND2_X1 U773 ( .A1(G2067), .A2(n940), .ZN(n688) );
  XNOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n691) );
  INV_X1 U775 ( .A(n691), .ZN(n686) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n686), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n689), .A2(n706), .ZN(n697) );
  INV_X1 U779 ( .A(G1341), .ZN(n946) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n940), .ZN(n951) );
  NAND2_X1 U781 ( .A1(n946), .A2(n951), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n722), .A2(n690), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n706), .A2(G1996), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n945), .A2(n695), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U789 ( .A1(G299), .A2(n700), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT28), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n705) );
  XOR2_X1 U792 ( .A(KEYINPUT95), .B(KEYINPUT29), .Z(n704) );
  XNOR2_X1 U793 ( .A(n705), .B(n704), .ZN(n710) );
  XOR2_X1 U794 ( .A(G2078), .B(KEYINPUT25), .Z(n917) );
  NOR2_X1 U795 ( .A1(n917), .A2(n722), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n706), .A2(G1961), .ZN(n707) );
  NOR2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n715) );
  NOR2_X1 U798 ( .A1(G301), .A2(n715), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n721) );
  NOR2_X1 U800 ( .A1(G1966), .A2(n761), .ZN(n736) );
  NOR2_X1 U801 ( .A1(G2084), .A2(n711), .ZN(n733) );
  NOR2_X1 U802 ( .A1(n736), .A2(n733), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G8), .A2(n712), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n713), .B(KEYINPUT30), .ZN(n714) );
  NOR2_X1 U805 ( .A1(G168), .A2(n714), .ZN(n717) );
  AND2_X1 U806 ( .A1(G301), .A2(n715), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U808 ( .A(n718), .B(KEYINPUT31), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT96), .B(n719), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n734), .A2(G286), .ZN(n729) );
  INV_X1 U811 ( .A(G8), .ZN(n727) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n761), .ZN(n724) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n722), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n725), .A2(G303), .ZN(n726) );
  OR2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U817 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n730) );
  NAND2_X1 U818 ( .A1(n733), .A2(G8), .ZN(n738) );
  INV_X1 U819 ( .A(n734), .ZN(n735) );
  NOR2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n738), .A2(n737), .ZN(n754) );
  NAND2_X1 U822 ( .A1(G288), .A2(G1976), .ZN(n739) );
  XOR2_X1 U823 ( .A(KEYINPUT99), .B(n739), .Z(n938) );
  AND2_X1 U824 ( .A1(n754), .A2(n938), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n753), .A2(n740), .ZN(n744) );
  INV_X1 U826 ( .A(n938), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n747) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U829 ( .A1(n747), .A2(n741), .ZN(n939) );
  OR2_X1 U830 ( .A1(n742), .A2(n939), .ZN(n743) );
  AND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n761), .A2(n745), .ZN(n746) );
  OR2_X1 U833 ( .A1(n746), .A2(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U834 ( .A1(n747), .A2(KEYINPUT33), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n748), .A2(n761), .ZN(n750) );
  XOR2_X1 U836 ( .A(G1981), .B(G305), .Z(n955) );
  INV_X1 U837 ( .A(n955), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U841 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U844 ( .A1(n758), .A2(n761), .ZN(n764) );
  NOR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U846 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  NOR2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U848 ( .A(n762), .B(KEYINPUT92), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n765) );
  AND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n799) );
  NAND2_X1 U851 ( .A1(n884), .A2(G140), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G104), .A2(n885), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT34), .B(n769), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G128), .A2(n891), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G116), .A2(n889), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U858 ( .A(n772), .B(KEYINPUT35), .Z(n773) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U860 ( .A(KEYINPUT36), .B(n775), .Z(n776) );
  XOR2_X1 U861 ( .A(KEYINPUT86), .B(n776), .Z(n871) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n802) );
  NOR2_X1 U863 ( .A1(n871), .A2(n802), .ZN(n979) );
  NAND2_X1 U864 ( .A1(n812), .A2(n979), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT87), .B(n777), .Z(n809) );
  INV_X1 U866 ( .A(n809), .ZN(n796) );
  NAND2_X1 U867 ( .A1(n891), .A2(G119), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G95), .A2(n885), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G131), .A2(n884), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G107), .A2(n889), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n866) );
  INV_X1 U874 ( .A(G1991), .ZN(n803) );
  NOR2_X1 U875 ( .A1(n866), .A2(n803), .ZN(n793) );
  NAND2_X1 U876 ( .A1(n885), .A2(G105), .ZN(n784) );
  XNOR2_X1 U877 ( .A(n784), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G141), .A2(n884), .ZN(n786) );
  NAND2_X1 U879 ( .A1(G129), .A2(n891), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n889), .A2(G117), .ZN(n787) );
  XOR2_X1 U882 ( .A(KEYINPUT88), .B(n787), .Z(n788) );
  NOR2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n870) );
  AND2_X1 U885 ( .A1(n870), .A2(G1996), .ZN(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n981) );
  INV_X1 U887 ( .A(n812), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n981), .A2(n794), .ZN(n806) );
  XOR2_X1 U889 ( .A(KEYINPUT89), .B(n806), .Z(n795) );
  NOR2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(n797), .Z(n798) );
  NOR2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n815) );
  NAND2_X1 U894 ( .A1(n871), .A2(n802), .ZN(n983) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n870), .ZN(n974) );
  AND2_X1 U896 ( .A1(n803), .A2(n866), .ZN(n968) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n968), .A2(n804), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n974), .A2(n807), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n983), .A2(n811), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U909 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n819) );
  XOR2_X1 U911 ( .A(KEYINPUT101), .B(n819), .Z(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(G188) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  INV_X1 U916 ( .A(G69), .ZN(G235) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U919 ( .A(G1348), .B(G2454), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n824), .B(G2430), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(G1341), .ZN(n831) );
  XOR2_X1 U922 ( .A(G2443), .B(G2427), .Z(n827) );
  XNOR2_X1 U923 ( .A(G2438), .B(G2446), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(n829) );
  XOR2_X1 U925 ( .A(G2451), .B(G2435), .Z(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n832), .A2(G14), .ZN(n833) );
  XOR2_X1 U929 ( .A(KEYINPUT100), .B(n833), .Z(G401) );
  XOR2_X1 U930 ( .A(G2100), .B(G2096), .Z(n835) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2072), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2084), .B(G2078), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1961), .B(G1966), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1981), .B(G1976), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G1971), .B(G1986), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT103), .B(G2474), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1956), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT102), .B(n852), .Z(G319) );
  NAND2_X1 U951 ( .A1(n884), .A2(G136), .ZN(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT104), .B(n853), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n891), .A2(G124), .ZN(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT44), .B(n854), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(KEYINPUT105), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G112), .A2(n889), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n885), .A2(G100), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT106), .B(n860), .Z(n861) );
  NOR2_X1 U961 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT111), .B(KEYINPUT108), .Z(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n865), .B(G162), .Z(n868) );
  XNOR2_X1 U966 ( .A(G160), .B(n866), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n869), .B(n967), .Z(n873) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n883) );
  NAND2_X1 U971 ( .A1(G130), .A2(n891), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G118), .A2(n889), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U974 ( .A1(G106), .A2(n885), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT107), .B(n876), .Z(n878) );
  NAND2_X1 U976 ( .A1(n884), .A2(G142), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(n879), .B(KEYINPUT45), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(n883), .B(n882), .Z(n898) );
  NAND2_X1 U981 ( .A1(n884), .A2(G139), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G103), .A2(n885), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(KEYINPUT109), .B(n888), .Z(n896) );
  NAND2_X1 U985 ( .A1(n889), .A2(G115), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n890), .B(KEYINPUT110), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G127), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n985) );
  XOR2_X1 U991 ( .A(n985), .B(G164), .Z(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U994 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n903) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U997 ( .A(G171), .B(G286), .Z(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1001 ( .A(KEYINPUT49), .B(n907), .Z(n908) );
  NAND2_X1 U1002 ( .A1(n908), .A2(G319), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n909), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(KEYINPUT114), .B(n910), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1009 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n992) );
  XOR2_X1 U1010 ( .A(G34), .B(KEYINPUT122), .Z(n914) );
  XNOR2_X1 U1011 ( .A(G2084), .B(KEYINPUT54), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n932) );
  XNOR2_X1 U1013 ( .A(G2090), .B(G35), .ZN(n930) );
  XNOR2_X1 U1014 ( .A(G25), .B(G1991), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n915), .B(KEYINPUT119), .ZN(n922) );
  XOR2_X1 U1016 ( .A(G32), .B(G1996), .Z(n916) );
  NAND2_X1 U1017 ( .A1(n916), .A2(G28), .ZN(n920) );
  XOR2_X1 U1018 ( .A(G27), .B(n917), .Z(n918) );
  XNOR2_X1 U1019 ( .A(KEYINPUT121), .B(n918), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G26), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G2072), .B(G33), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1025 ( .A(KEYINPUT120), .B(n925), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n992), .B(n933), .ZN(n935) );
  INV_X1 U1031 ( .A(G29), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(G11), .A2(n936), .ZN(n966) );
  XNOR2_X1 U1034 ( .A(G16), .B(KEYINPUT123), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(n937), .B(KEYINPUT56), .ZN(n963) );
  XNOR2_X1 U1036 ( .A(G1961), .B(G171), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(G1348), .A2(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n961) );
  XNOR2_X1 U1041 ( .A(n946), .B(n945), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(G1971), .A2(G303), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(G1956), .B(G299), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(G168), .B(G1966), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT57), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n964), .B(KEYINPUT124), .ZN(n965) );
  NOR2_X1 U1055 ( .A1(n966), .A2(n965), .ZN(n996) );
  XOR2_X1 U1056 ( .A(G160), .B(G2084), .Z(n971) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT115), .B(n969), .ZN(n970) );
  NOR2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1060 ( .A(KEYINPUT116), .B(n972), .ZN(n977) );
  XOR2_X1 U1061 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1063 ( .A(KEYINPUT51), .B(n975), .Z(n976) );
  NAND2_X1 U1064 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1065 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1066 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1067 ( .A(n982), .B(KEYINPUT117), .ZN(n984) );
  NAND2_X1 U1068 ( .A1(n984), .A2(n983), .ZN(n990) );
  XOR2_X1 U1069 ( .A(G2072), .B(n985), .Z(n987) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n986) );
  NOR2_X1 U1071 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1072 ( .A(KEYINPUT50), .B(n988), .Z(n989) );
  NOR2_X1 U1073 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1074 ( .A(KEYINPUT52), .B(n991), .ZN(n993) );
  NAND2_X1 U1075 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1076 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1077 ( .A1(n996), .A2(n995), .ZN(n1022) );
  XOR2_X1 U1078 ( .A(G1986), .B(G24), .Z(n1000) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n998) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n997) );
  NOR2_X1 U1081 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1082 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1083 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(n1002), .B(n1001), .ZN(n1015) );
  XNOR2_X1 U1085 ( .A(KEYINPUT59), .B(G1348), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(n1003), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n1008) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(G19), .B(G1341), .ZN(n1004) );
  NOR2_X1 U1090 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1092 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G5), .ZN(n1012) );
  NOR2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1097 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1098 ( .A(G21), .B(G1966), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1100 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NOR2_X1 U1102 ( .A1(G16), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1103 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1104 ( .A(n1023), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

