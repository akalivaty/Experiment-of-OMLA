//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT73), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT72), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(G125), .A2(G140), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n190), .B(KEYINPUT16), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n197), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n187), .B2(new_n191), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n190), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n193), .A2(new_n195), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n197), .B1(new_n206), .B2(G140), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT73), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n198), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(G146), .A3(new_n189), .ZN(new_n211));
  OR2_X1    g025(.A1(KEYINPUT88), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT88), .A2(G143), .ZN(new_n213));
  NOR2_X1   g027(.A1(G237), .A2(G953), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(G214), .ZN(new_n215));
  INV_X1    g029(.A(G237), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G214), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT88), .A2(G143), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n213), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n218), .B1(new_n224), .B2(new_n219), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n212), .A2(G214), .A3(new_n214), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n223), .B1(new_n230), .B2(new_n222), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n205), .A2(new_n211), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n227), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(new_n233), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(G146), .B(new_n200), .C1(new_n187), .C2(new_n191), .ZN(new_n239));
  XNOR2_X1  g053(.A(G125), .B(G140), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n204), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT90), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n238), .A2(new_n244), .A3(KEYINPUT91), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n221), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n236), .B1(new_n248), .B2(new_n233), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n239), .A2(new_n241), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n239), .A2(KEYINPUT90), .A3(new_n241), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n232), .B1(new_n245), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G113), .B(G122), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT92), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(G104), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT91), .B1(new_n238), .B2(new_n244), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n249), .A2(new_n254), .A3(new_n246), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT19), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n240), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n201), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n230), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n259), .B1(new_n267), .B2(new_n211), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n256), .A2(new_n259), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n270));
  NOR2_X1   g084(.A1(G475), .A2(G902), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n269), .A2(KEYINPUT93), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n262), .A2(new_n268), .ZN(new_n275));
  AOI21_X1  g089(.A(G146), .B1(new_n210), .B2(new_n189), .ZN(new_n276));
  AOI211_X1 g090(.A(new_n204), .B(new_n188), .C1(new_n209), .C2(new_n198), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n231), .B1(new_n260), .B2(new_n261), .ZN(new_n279));
  INV_X1    g093(.A(new_n259), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n274), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(KEYINPUT94), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n256), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  INV_X1    g099(.A(new_n283), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n262), .A3(new_n232), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n284), .A2(KEYINPUT95), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G475), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n256), .B2(new_n283), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT95), .B1(new_n290), .B2(new_n287), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n273), .A2(new_n282), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT14), .A3(G122), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G122), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(G107), .B(new_n295), .C1(new_n297), .C2(KEYINPUT14), .ZN(new_n298));
  INV_X1    g112(.A(G107), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(G128), .B(G143), .Z(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT67), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G134), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n301), .A2(new_n306), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n298), .B(new_n300), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n296), .B(G107), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT13), .ZN(new_n311));
  INV_X1    g125(.A(G143), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G128), .ZN(new_n313));
  OAI211_X1 g127(.A(G134), .B(new_n313), .C1(new_n301), .C2(new_n311), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n306), .B2(new_n301), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT9), .B(G234), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n317), .A2(new_n318), .A3(G953), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n316), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n285), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT15), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G478), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(G478), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n285), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G952), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(G234), .A2(G237), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(G902), .A3(G953), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT21), .B(G898), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G221), .B1(new_n317), .B2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n299), .A2(G104), .ZN(new_n340));
  INV_X1    g154(.A(G104), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G107), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(KEYINPUT3), .A3(G107), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n299), .A2(G104), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n341), .B2(G107), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(KEYINPUT76), .A3(new_n339), .A4(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n299), .A3(G104), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n350), .A3(new_n339), .A4(new_n342), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n204), .A3(G143), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n312), .A2(G146), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT66), .B1(new_n312), .B2(G146), .ZN(new_n360));
  INV_X1    g174(.A(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT1), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n356), .A3(new_n357), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(G143), .B2(new_n204), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n360), .A2(new_n356), .A3(new_n357), .A4(new_n362), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n354), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n347), .A2(new_n350), .A3(new_n342), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n351), .A2(new_n352), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n351), .A2(new_n352), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT4), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT0), .A2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G143), .B(G146), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT65), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n204), .A2(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n357), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n380), .A4(new_n379), .ZN(new_n387));
  INV_X1    g201(.A(new_n380), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n360), .A2(new_n356), .A3(new_n388), .A4(new_n357), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n374), .A2(G101), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT78), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n374), .A2(new_n392), .A3(new_n395), .A4(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n378), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT11), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n399), .A2(new_n302), .A3(G137), .ZN(new_n400));
  AOI21_X1  g214(.A(G137), .B1(new_n303), .B2(new_n305), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n402), .B2(new_n399), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT67), .B(G134), .ZN(new_n404));
  AOI21_X1  g218(.A(G131), .B1(new_n404), .B2(G137), .ZN(new_n405));
  INV_X1    g219(.A(new_n400), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n303), .A2(new_n305), .A3(G137), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n406), .B(new_n407), .C1(new_n401), .C2(KEYINPUT11), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n403), .A2(new_n405), .B1(new_n408), .B2(G131), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n385), .B1(new_n366), .B2(new_n361), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n368), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n354), .A2(KEYINPUT10), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n373), .A2(new_n398), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(G227), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n414), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT12), .ZN(new_n420));
  INV_X1    g234(.A(new_n343), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n376), .B2(new_n377), .ZN(new_n422));
  INV_X1    g236(.A(new_n411), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n420), .B(new_n409), .C1(new_n424), .C2(new_n371), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n409), .B1(new_n424), .B2(new_n371), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(KEYINPUT12), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n419), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n373), .A2(new_n398), .A3(new_n412), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n408), .A2(G131), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n399), .B1(new_n404), .B2(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n405), .A3(new_n406), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n413), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n417), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT80), .B(G469), .Z(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n285), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n413), .B1(new_n427), .B2(new_n425), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n441), .A2(new_n417), .B1(new_n419), .B2(new_n434), .ZN(new_n442));
  OAI21_X1  g256(.A(G469), .B1(new_n442), .B2(G902), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n338), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n293), .A2(new_n336), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G214), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n390), .A2(new_n447), .A3(new_n206), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n390), .B2(new_n206), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n411), .A2(new_n206), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G224), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT7), .B1(new_n452), .B2(G953), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n451), .A2(KEYINPUT85), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n390), .A2(new_n206), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n457), .B2(KEYINPUT82), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n390), .A2(new_n447), .A3(new_n206), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n460), .B2(new_n453), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT84), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT8), .Z(new_n465));
  XNOR2_X1  g279(.A(G116), .B(G119), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n294), .A2(KEYINPUT5), .ZN(new_n469));
  INV_X1    g283(.A(G119), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT2), .B(G113), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n467), .A2(new_n471), .B1(new_n473), .B2(new_n466), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n354), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n354), .A2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n465), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n472), .B(new_n466), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n394), .B2(new_n396), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n378), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n475), .A3(new_n463), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n458), .A2(new_n459), .A3(new_n454), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n462), .B2(new_n485), .ZN(new_n486));
  NOR4_X1   g300(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT83), .A4(new_n450), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n458), .B2(new_n459), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n487), .A2(new_n489), .B1(new_n452), .B2(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n452), .A2(G953), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n458), .A2(new_n488), .A3(new_n459), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n480), .A2(new_n378), .B1(new_n354), .B2(new_n474), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n463), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n496), .B2(new_n463), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n496), .A2(new_n463), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n486), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n486), .A2(new_n506), .A3(new_n510), .A4(new_n507), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n507), .B(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n497), .A2(new_n498), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n482), .A2(new_n500), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n515), .A2(new_n501), .B1(new_n490), .B2(new_n494), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT85), .B1(new_n451), .B2(new_n454), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n460), .A2(new_n456), .A3(new_n453), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n285), .B1(new_n519), .B2(new_n484), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n512), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n446), .B1(new_n509), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n445), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT75), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT22), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(G137), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n361), .A2(G119), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n470), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G110), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n361), .A2(KEYINPUT23), .A3(G119), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n470), .A2(G128), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n533), .C1(new_n538), .C2(KEYINPUT23), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(G110), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n205), .B2(new_n211), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n534), .A2(new_n535), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n539), .B2(G110), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n241), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n548), .A2(new_n211), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n531), .B1(new_n542), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n540), .B1(new_n276), .B2(new_n277), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n211), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n530), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n527), .B1(new_n554), .B2(G902), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n285), .A3(new_n553), .A4(new_n526), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n318), .B1(G234), .B2(new_n285), .ZN(new_n558));
  INV_X1    g372(.A(new_n554), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(G902), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n557), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G137), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G134), .ZN(new_n563));
  OAI21_X1  g377(.A(G131), .B1(new_n401), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n432), .A2(new_n411), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n479), .C1(new_n409), .C2(new_n390), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT28), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n479), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n390), .B1(new_n430), .B2(new_n432), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n432), .A2(new_n411), .A3(new_n564), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(new_n566), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT27), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n214), .A2(new_n576), .A3(G210), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n214), .B2(G210), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT26), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n579), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT26), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n577), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n580), .A2(new_n583), .A3(G101), .ZN(new_n584));
  AOI21_X1  g398(.A(G101), .B1(new_n580), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n575), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(KEYINPUT70), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT70), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n573), .A2(new_n596), .A3(new_n566), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT71), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT28), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n595), .B(new_n568), .C1(new_n597), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n588), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n602));
  NAND2_X1  g416(.A1(new_n433), .A2(new_n391), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n565), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n565), .A2(KEYINPUT30), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n570), .B1(new_n605), .B2(new_n571), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT68), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n602), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n571), .B2(new_n572), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT30), .B(new_n565), .C1(new_n409), .C2(new_n390), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT68), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n570), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n586), .B1(new_n613), .B2(new_n566), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n590), .B1(new_n601), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  NOR2_X1   g430(.A1(G472), .A2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n566), .A2(new_n586), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n607), .B2(new_n612), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT31), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n598), .A2(KEYINPUT28), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n573), .A2(new_n596), .A3(new_n566), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n569), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI22_X1  g437(.A1(new_n619), .A2(new_n620), .B1(new_n623), .B2(new_n595), .ZN(new_n624));
  INV_X1    g438(.A(new_n618), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n613), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(KEYINPUT32), .B(new_n617), .C1(new_n624), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n616), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n568), .B1(new_n597), .B2(new_n599), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n594), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n632), .B(new_n627), .C1(new_n620), .C2(new_n619), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT32), .B1(new_n633), .B2(new_n617), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n561), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n524), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT96), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  AND2_X1   g453(.A1(new_n633), .A2(new_n617), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n633), .B2(new_n285), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(KEYINPUT97), .A3(new_n561), .A4(new_n444), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n444), .A2(new_n561), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n633), .A2(new_n617), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n613), .A2(new_n625), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n648), .A2(KEYINPUT31), .B1(new_n594), .B2(new_n631), .ZN(new_n649));
  AOI21_X1  g463(.A(G902), .B1(new_n649), .B2(new_n627), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n647), .B1(new_n650), .B2(new_n641), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n645), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n320), .B(KEYINPUT33), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n285), .A2(G478), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT98), .B(G478), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n654), .A2(new_n656), .B1(new_n321), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n281), .A2(new_n270), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n275), .B(new_n271), .C1(new_n279), .C2(new_n280), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n272), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT95), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n285), .B1(new_n279), .B2(new_n286), .ZN(new_n664));
  INV_X1    g478(.A(new_n287), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(G475), .A3(new_n288), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n658), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n335), .ZN(new_n670));
  INV_X1    g484(.A(new_n446), .ZN(new_n671));
  INV_X1    g485(.A(new_n507), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n516), .B2(new_n520), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n671), .B1(new_n673), .B2(new_n508), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n653), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT34), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n341), .ZN(G6));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n508), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n446), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n660), .A2(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n667), .A2(new_n326), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n335), .B(KEYINPUT99), .Z(new_n685));
  NAND3_X1  g499(.A1(new_n653), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT35), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n299), .ZN(G9));
  NAND2_X1  g502(.A1(new_n557), .A2(new_n558), .ZN(new_n689));
  OAI22_X1  g503(.A1(new_n542), .A2(new_n549), .B1(KEYINPUT36), .B2(new_n531), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n531), .A2(KEYINPUT36), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n551), .A2(new_n552), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n560), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n651), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n524), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(G900), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n333), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n330), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n667), .A2(new_n682), .A3(new_n326), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n630), .B2(new_n634), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n444), .A3(new_n674), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n695), .A2(new_n444), .A3(new_n674), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT32), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n647), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n629), .A3(new_n616), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(KEYINPUT101), .A3(new_n712), .A4(new_n705), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  NAND2_X1  g529(.A1(new_n573), .A2(new_n566), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n594), .A3(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n594), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n648), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n641), .B1(new_n721), .B2(new_n285), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n647), .B2(new_n710), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(KEYINPUT103), .A3(new_n629), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT103), .B1(new_n723), .B2(new_n629), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n695), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n511), .A2(new_n521), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT38), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT38), .B1(new_n509), .B2(new_n522), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n704), .B(KEYINPUT39), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n444), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT40), .Z(new_n736));
  AOI22_X1  g550(.A1(new_n662), .A2(new_n667), .B1(new_n323), .B2(new_n325), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(new_n446), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n727), .A2(new_n733), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  INV_X1    g554(.A(new_n658), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n292), .A2(new_n741), .A3(new_n704), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n709), .A2(new_n743), .A3(new_n712), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  INV_X1    g559(.A(G469), .ZN(new_n746));
  AOI21_X1  g560(.A(G902), .B1(new_n428), .B2(new_n436), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n440), .B(new_n337), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n679), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n636), .A2(new_n670), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT41), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G113), .ZN(G15));
  INV_X1    g566(.A(new_n685), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n636), .A2(new_n684), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G116), .ZN(G18));
  NOR3_X1   g570(.A1(new_n696), .A2(new_n679), .A3(new_n748), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n292), .A2(new_n335), .A3(new_n326), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n712), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND3_X1  g574(.A1(new_n674), .A2(new_n292), .A3(new_n326), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n763));
  OAI22_X1  g577(.A1(new_n619), .A2(new_n620), .B1(new_n575), .B2(new_n595), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n628), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n642), .B1(new_n766), .B2(new_n617), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n762), .A2(new_n767), .A3(new_n561), .A4(new_n754), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND2_X1  g583(.A1(new_n742), .A2(KEYINPUT105), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n668), .A2(new_n771), .A3(new_n704), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n757), .A2(new_n767), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  NAND4_X1  g588(.A1(new_n730), .A2(new_n446), .A3(new_n521), .A4(new_n511), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n434), .A2(new_n413), .A3(new_n418), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n354), .A2(new_n370), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n354), .A2(new_n411), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n433), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n420), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n426), .A2(KEYINPUT12), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n373), .A2(new_n398), .A3(new_n412), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n409), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n776), .B1(new_n783), .B2(new_n418), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n746), .B1(new_n784), .B2(new_n285), .ZN(new_n785));
  AOI211_X1 g599(.A(G902), .B(new_n438), .C1(new_n428), .C2(new_n436), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n337), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n770), .A2(new_n772), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n629), .B(new_n616), .C1(new_n634), .C2(KEYINPUT106), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n634), .A2(KEYINPUT106), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n561), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT42), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n444), .A2(new_n728), .A3(new_n446), .A4(new_n730), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n635), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n770), .A4(new_n772), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT107), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n226), .ZN(G33));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n705), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NOR2_X1   g616(.A1(new_n746), .A2(new_n285), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT45), .B(new_n776), .C1(new_n783), .C2(new_n418), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n442), .A2(new_n806), .A3(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(G469), .B1(new_n442), .B2(KEYINPUT45), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n803), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n440), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n809), .B1(new_n805), .B2(new_n807), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT46), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(new_n803), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n337), .B(new_n734), .C1(new_n812), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n813), .B2(new_n803), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(new_n440), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT109), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n337), .A4(new_n734), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT43), .B1(new_n292), .B2(new_n658), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT43), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n662), .A2(new_n741), .A3(new_n824), .A4(new_n667), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n651), .A3(new_n695), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n775), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n817), .A2(new_n822), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  NAND2_X1  g645(.A1(new_n820), .A2(new_n337), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT47), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n712), .A2(new_n742), .A3(new_n561), .A4(new_n775), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT47), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n820), .A2(new_n835), .A3(new_n337), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  NAND2_X1  g652(.A1(new_n327), .A2(new_n217), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n326), .B(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n293), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n523), .B1(new_n841), .B2(new_n669), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n652), .A3(new_n644), .A4(new_n685), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n524), .B1(new_n636), .B2(new_n697), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n788), .A2(new_n695), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n770), .A2(new_n772), .A3(new_n767), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n840), .B1(new_n330), .B2(new_n703), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n712), .A2(new_n848), .A3(new_n667), .A4(new_n682), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n636), .A2(new_n705), .A3(new_n788), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n845), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n750), .A2(new_n755), .A3(new_n768), .A4(new_n759), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n798), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n762), .A2(new_n754), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n767), .A2(new_n561), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n749), .A2(new_n695), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n712), .A2(new_n758), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n857), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n335), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n749), .A2(new_n862), .A3(new_n668), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n684), .A2(new_n754), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n635), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n793), .A4(new_n797), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n853), .A2(new_n856), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n444), .A2(new_n704), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n761), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n696), .B(new_n870), .C1(new_n724), .C2(new_n725), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(KEYINPUT52), .A3(new_n744), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n714), .A2(new_n873), .A3(new_n773), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n714), .B2(new_n773), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n714), .A2(new_n871), .A3(new_n744), .A4(new_n773), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n877), .A2(KEYINPUT113), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT113), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n868), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n877), .B(KEYINPUT52), .ZN(new_n884));
  INV_X1    g698(.A(new_n798), .ZN(new_n885));
  INV_X1    g699(.A(new_n845), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n850), .A2(new_n852), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n866), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n851), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n881), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT53), .B1(new_n884), .B2(new_n888), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(KEYINPUT54), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n747), .A2(new_n746), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n786), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n833), .A2(new_n836), .B1(new_n338), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n338), .ZN(new_n900));
  INV_X1    g714(.A(new_n836), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n835), .B1(new_n820), .B2(new_n337), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n775), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n823), .A2(new_n331), .A3(new_n825), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(KEYINPUT115), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT115), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n858), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n899), .A2(new_n905), .A3(new_n906), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n907), .B(KEYINPUT115), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n775), .A2(new_n748), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT118), .Z(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n914), .A3(new_n695), .A4(new_n767), .ZN(new_n915));
  INV_X1    g729(.A(new_n561), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n330), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n292), .A2(new_n741), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n914), .A2(new_n726), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n915), .A2(KEYINPUT51), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n733), .A2(new_n446), .A3(new_n748), .ZN(new_n923));
  INV_X1    g737(.A(new_n858), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n912), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT116), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT116), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n910), .A2(new_n927), .A3(new_n923), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n922), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n910), .A2(KEYINPUT50), .A3(new_n923), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n911), .B(new_n920), .C1(new_n929), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n910), .A2(new_n749), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n914), .A2(new_n668), .A3(new_n726), .A4(new_n917), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n934), .A3(new_n328), .ZN(new_n935));
  INV_X1    g749(.A(new_n792), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n912), .A2(new_n914), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT48), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n910), .A2(new_n906), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n919), .B(new_n915), .C1(new_n941), .C2(new_n898), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n926), .A2(new_n928), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n921), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n932), .B(new_n940), .C1(new_n945), .C2(KEYINPUT51), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n839), .B1(new_n895), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n561), .A2(new_n446), .A3(new_n337), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n948), .A2(new_n292), .A3(new_n658), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT110), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n897), .B(KEYINPUT49), .Z(new_n953));
  NOR4_X1   g767(.A1(new_n951), .A2(new_n952), .A3(new_n733), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n726), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n947), .A2(KEYINPUT120), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G75));
  NOR2_X1   g774(.A1(new_n217), .A2(G952), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT121), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n285), .B1(new_n882), .B2(new_n889), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n512), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n495), .A2(new_n505), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n516), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT56), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n963), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT56), .B1(new_n964), .B2(G210), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n972), .B(KEYINPUT122), .C1(new_n968), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n964), .A2(G210), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n968), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  INV_X1    g791(.A(new_n512), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n285), .B(new_n978), .C1(new_n882), .C2(new_n889), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n962), .B1(new_n979), .B2(new_n970), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n974), .A2(new_n981), .ZN(G51));
  NAND3_X1  g796(.A1(new_n853), .A2(new_n856), .A3(new_n867), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n877), .A2(new_n878), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n877), .A2(KEYINPUT113), .A3(new_n878), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n988), .B2(new_n876), .ZN(new_n989));
  INV_X1    g803(.A(new_n888), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n877), .B(new_n878), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT53), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT54), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(KEYINPUT123), .A3(new_n890), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n882), .A2(new_n889), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT54), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n803), .B(KEYINPUT57), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n437), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n964), .A2(new_n813), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n961), .B1(new_n1000), .B2(new_n1001), .ZN(G54));
  NAND2_X1  g816(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n964), .A2(new_n269), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n269), .B1(new_n964), .B2(new_n1004), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n961), .ZN(G60));
  NAND2_X1  g821(.A1(G478), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT59), .Z(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n890), .B2(new_n894), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n962), .B1(new_n1010), .B2(new_n654), .ZN(new_n1011));
  INV_X1    g825(.A(new_n654), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(new_n1009), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n994), .A2(new_n997), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT124), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n994), .A2(new_n1016), .A3(new_n997), .A4(new_n1013), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1011), .B1(new_n1015), .B2(new_n1017), .ZN(G63));
  NOR2_X1   g832(.A1(new_n989), .A2(new_n992), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G217), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT60), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n554), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1021), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n995), .A2(new_n692), .A3(new_n690), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1022), .A2(new_n962), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT61), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(G66));
  NAND2_X1  g841(.A1(new_n886), .A2(new_n866), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G224), .A2(G953), .ZN(new_n1029));
  OAI22_X1  g843(.A1(new_n1028), .A2(G953), .B1(new_n334), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n515), .B(new_n501), .C1(G898), .C2(new_n217), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1030), .B(new_n1031), .Z(G69));
  OAI21_X1  g846(.A(G953), .B1(new_n415), .B2(new_n702), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1033), .B(KEYINPUT127), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n609), .A2(new_n610), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(new_n265), .Z(new_n1037));
  NAND2_X1  g851(.A1(new_n702), .A2(G953), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n744), .B1(new_n874), .B2(new_n875), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n793), .A2(new_n797), .A3(new_n801), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n817), .A2(new_n762), .A3(new_n936), .A4(new_n822), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n830), .A2(new_n837), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1038), .B1(new_n1044), .B2(G953), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1037), .B1(new_n1045), .B2(KEYINPUT126), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n1047), .B(new_n1038), .C1(new_n1044), .C2(G953), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n739), .B(new_n744), .C1(new_n874), .C2(new_n875), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT62), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n714), .A2(new_n773), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n714), .A2(new_n873), .A3(new_n773), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1055), .A2(KEYINPUT62), .A3(new_n739), .A4(new_n744), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n841), .A2(new_n669), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n795), .A2(new_n734), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n830), .A2(new_n837), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(KEYINPUT125), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT125), .ZN(new_n1063));
  AOI211_X1 g877(.A(new_n1063), .B(new_n1060), .C1(new_n1051), .C2(new_n1056), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n217), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI221_X4 g879(.A(new_n1035), .B1(new_n1046), .B2(new_n1048), .C1(new_n1065), .C2(new_n1037), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1065), .A2(new_n1037), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1034), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g883(.A1(new_n1066), .A2(new_n1069), .ZN(G72));
  NAND3_X1  g884(.A1(new_n1044), .A2(new_n866), .A3(new_n886), .ZN(new_n1071));
  NAND2_X1  g885(.A1(G472), .A2(G902), .ZN(new_n1072));
  XOR2_X1   g886(.A(new_n1072), .B(KEYINPUT63), .Z(new_n1073));
  NAND2_X1  g887(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g888(.A1(new_n1074), .A2(new_n613), .A3(new_n587), .A4(new_n566), .ZN(new_n1075));
  INV_X1    g889(.A(new_n961), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n892), .A2(new_n893), .ZN(new_n1077));
  OAI21_X1  g891(.A(new_n1073), .B1(new_n614), .B2(new_n619), .ZN(new_n1078));
  OAI211_X1 g892(.A(new_n1075), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  OR2_X1    g893(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1080));
  OAI21_X1  g894(.A(new_n1073), .B1(new_n1080), .B2(new_n1028), .ZN(new_n1081));
  AOI21_X1  g895(.A(new_n587), .B1(new_n613), .B2(new_n566), .ZN(new_n1082));
  AOI21_X1  g896(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(G57));
endmodule


