//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT80), .B(G469), .Z(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(G101), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT75), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT75), .A4(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n213), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G143), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G101), .B1(new_n198), .B2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n199), .A2(new_n221), .A3(new_n202), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n204), .A2(G101), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n201), .A2(G104), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n198), .A2(G107), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n222), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n232));
  OAI211_X1 g046(.A(G128), .B(new_n232), .C1(new_n216), .C2(new_n217), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n212), .B(new_n214), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT10), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n231), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n226), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n229), .A2(new_n222), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n235), .A4(new_n233), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n233), .A2(new_n229), .A3(new_n222), .A4(new_n235), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT76), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n248), .B2(new_n237), .ZN(new_n249));
  AOI211_X1 g063(.A(KEYINPUT77), .B(KEYINPUT10), .C1(new_n245), .C2(new_n247), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n241), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT79), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G131), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n258), .A3(new_n262), .A4(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT79), .B(new_n241), .C1(new_n249), .C2(new_n250), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n253), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n264), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n267), .B(new_n241), .C1(new_n249), .C2(new_n250), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n197), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n197), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n246), .B(new_n244), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n233), .A2(new_n235), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n243), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT12), .B(new_n264), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n245), .B2(new_n247), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n267), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n270), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n190), .B(new_n192), .C1(new_n269), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n274), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n197), .B1(new_n268), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n226), .A2(new_n240), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT77), .B1(new_n271), .B2(KEYINPUT10), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n248), .A2(new_n242), .A3(new_n237), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n196), .B1(new_n285), .B2(new_n267), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n266), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G469), .B1(new_n287), .B2(G902), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n191), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G475), .A2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G143), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n213), .A2(KEYINPUT88), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G237), .A2(G953), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G214), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(G214), .A3(new_n296), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT18), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(new_n262), .ZN(new_n301));
  XNOR2_X1  g115(.A(G125), .B(G140), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(new_n211), .ZN(new_n303));
  INV_X1    g117(.A(new_n299), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(G214), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n301), .B(new_n303), .C1(new_n306), .C2(new_n300), .ZN(new_n307));
  XNOR2_X1  g121(.A(G113), .B(G122), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(new_n198), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n298), .A2(new_n262), .A3(new_n299), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT17), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n321), .A2(new_n313), .A3(new_n314), .A4(G125), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n211), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT17), .B(G131), .C1(new_n304), .C2(new_n305), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n316), .A2(new_n320), .A3(G146), .A4(new_n322), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n307), .B(new_n309), .C1(new_n312), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT90), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n324), .A3(new_n326), .A4(new_n325), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(KEYINPUT90), .A3(new_n309), .A4(new_n307), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n306), .A2(new_n310), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT89), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n306), .A2(new_n310), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n317), .A2(new_n319), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT19), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n302), .A2(KEYINPUT19), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n211), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n336), .A2(new_n326), .A3(new_n338), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n307), .ZN(new_n346));
  INV_X1    g160(.A(new_n309), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n291), .B1(new_n334), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n334), .A2(new_n348), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n354), .A2(KEYINPUT91), .A3(new_n350), .A4(new_n290), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n330), .A2(new_n333), .B1(new_n346), .B2(new_n347), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n356), .B2(new_n291), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n309), .B1(new_n332), .B2(new_n307), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n330), .B2(new_n333), .ZN(new_n360));
  OAI21_X1  g174(.A(G475), .B1(new_n360), .B2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n213), .A2(G128), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n234), .A2(G143), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G134), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n255), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  INV_X1    g183(.A(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G122), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n371), .A3(new_n201), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(KEYINPUT14), .A3(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n371), .ZN(new_n374));
  OAI211_X1 g188(.A(G107), .B(new_n373), .C1(new_n374), .C2(KEYINPUT14), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n367), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(G107), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n377), .A2(new_n372), .A3(KEYINPUT92), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT92), .B1(new_n377), .B2(new_n372), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n363), .B1(new_n362), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n362), .A2(new_n381), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT93), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT93), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n362), .A2(new_n385), .A3(new_n381), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n366), .B1(new_n387), .B2(new_n255), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n376), .B1(new_n380), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n188), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n376), .B(new_n391), .C1(new_n380), .C2(new_n388), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT94), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n190), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G478), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT95), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(G234), .A2(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G952), .A3(new_n194), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT21), .B(G898), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(G902), .A3(G953), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n404), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n395), .A2(new_n190), .A3(new_n397), .A4(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n405), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n358), .A2(new_n361), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n289), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G122), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G119), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G116), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n370), .A2(G119), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n223), .A2(new_n224), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT81), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n210), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n435));
  OAI21_X1  g249(.A(G113), .B1(new_n435), .B2(new_n425), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n435), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n434), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n231), .A3(new_n239), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n432), .B1(new_n431), .B2(new_n210), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n423), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n431), .A2(new_n210), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(new_n422), .A3(new_n441), .A4(new_n433), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n220), .B2(G125), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n220), .A2(new_n449), .A3(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n236), .A2(new_n318), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n194), .A2(G224), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT84), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n423), .C1(new_n442), .C2(new_n443), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n448), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n461), .A3(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n452), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n450), .ZN(new_n466));
  INV_X1    g280(.A(new_n463), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n466), .B(new_n453), .C1(new_n461), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT5), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(G113), .C1(new_n425), .C2(new_n435), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n243), .A2(new_n429), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n440), .B2(new_n243), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n422), .B(KEYINPUT8), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT85), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n476));
  INV_X1    g290(.A(new_n439), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n429), .B1(new_n477), .B2(new_n436), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n230), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n476), .B(new_n473), .C1(new_n479), .C2(new_n471), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n464), .B(new_n468), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n447), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n190), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n421), .B1(new_n460), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n483), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n448), .A2(new_n457), .A3(new_n459), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n420), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n419), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n417), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n424), .A2(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n234), .A2(G119), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT24), .B(G110), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT23), .A2(G119), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(G128), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n234), .A2(KEYINPUT66), .A3(KEYINPUT23), .A4(G119), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT67), .B(KEYINPUT23), .C1(new_n234), .C2(G119), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n494), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT67), .B1(new_n493), .B2(KEYINPUT23), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n497), .B1(new_n506), .B2(G110), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(new_n326), .C1(G146), .C2(new_n339), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n495), .A2(new_n496), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n324), .B2(new_n326), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(KEYINPUT68), .A3(G110), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT68), .B1(new_n506), .B2(G110), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n509), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n506), .A2(G110), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n509), .B1(new_n520), .B2(new_n511), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n508), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n508), .B(new_n525), .C1(new_n516), .C2(new_n521), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n190), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT71), .A4(new_n190), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n527), .A2(new_n190), .A3(new_n528), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT72), .B1(new_n535), .B2(KEYINPUT25), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n390), .B1(G234), .B2(new_n190), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n531), .A2(KEYINPUT72), .A3(new_n532), .A4(new_n533), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n527), .A2(new_n528), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n538), .A2(G902), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n296), .A2(G210), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT27), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n429), .A2(new_n430), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n257), .A2(G134), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n259), .A3(KEYINPUT64), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(G131), .C1(KEYINPUT64), .C2(new_n554), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n272), .A2(new_n263), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n220), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT65), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n558), .A2(new_n264), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n558), .B2(new_n264), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n553), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n264), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n557), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(KEYINPUT30), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n551), .B(new_n562), .C1(new_n568), .C2(new_n553), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT31), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n272), .A2(new_n263), .A3(new_n556), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(KEYINPUT65), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n558), .A2(new_n264), .A3(new_n559), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n565), .B1(new_n574), .B2(new_n564), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n552), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n551), .A4(new_n562), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n557), .A2(new_n563), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n552), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n552), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n581), .B(new_n582), .C1(new_n562), .C2(new_n579), .ZN(new_n583));
  INV_X1    g397(.A(new_n551), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n570), .A2(new_n578), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(KEYINPUT32), .A3(new_n587), .ZN(new_n591));
  INV_X1    g405(.A(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n567), .A2(new_n552), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n562), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n594), .B2(KEYINPUT28), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT29), .A3(new_n551), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n190), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT29), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n583), .B2(new_n584), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n576), .A2(new_n562), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n584), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n590), .A2(new_n591), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n547), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n460), .A2(new_n483), .A3(new_n421), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n420), .B1(new_n485), .B2(new_n486), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n418), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n489), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n289), .A3(new_n610), .A4(new_n416), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT96), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n492), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT97), .B(G101), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  NAND2_X1  g429(.A1(new_n586), .A2(new_n190), .ZN(new_n616));
  NAND2_X1  g430(.A1(KEYINPUT98), .A2(G472), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n546), .A2(new_n618), .A3(new_n540), .A4(new_n289), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n488), .A2(new_n411), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n355), .A2(new_n357), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT91), .B1(new_n349), .B2(new_n350), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n361), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n398), .A2(new_n399), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n395), .A2(new_n625), .A3(new_n397), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n393), .A2(KEYINPUT33), .A3(new_n394), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n393), .A2(new_n629), .A3(KEYINPUT33), .A4(new_n394), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n190), .A2(G478), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n620), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND2_X1  g452(.A1(new_n405), .A2(new_n413), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n351), .A2(new_n357), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n361), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n488), .A2(new_n411), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n619), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n522), .B(new_n647), .Z(new_n648));
  INV_X1    g462(.A(new_n545), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n539), .A2(new_n538), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT72), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n529), .B2(new_n532), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT25), .B1(new_n529), .B2(new_n530), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n533), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n646), .B(new_n651), .C1(new_n652), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n646), .B1(new_n540), .B2(new_n651), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n492), .A3(new_n612), .A4(new_n618), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AND3_X1   g477(.A1(new_n289), .A2(new_n603), .A3(new_n488), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n651), .B1(new_n652), .B2(new_n656), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n194), .A2(G900), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(G902), .A3(new_n406), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n407), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n640), .A2(new_n361), .A3(new_n639), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT102), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n664), .A2(new_n666), .A3(new_n657), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NAND2_X1  g489(.A1(new_n623), .A2(new_n639), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n418), .ZN(new_n678));
  OR3_X1    g492(.A1(new_n678), .A2(new_n665), .A3(KEYINPUT103), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT103), .B1(new_n678), .B2(new_n665), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n671), .B(KEYINPUT39), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n289), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n484), .A2(new_n487), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n289), .A2(new_n689), .A3(new_n682), .ZN(new_n690));
  INV_X1    g504(.A(G472), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n600), .A2(new_n551), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n594), .A2(new_n551), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(G902), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n590), .A2(new_n591), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n684), .A2(new_n688), .A3(new_n690), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n681), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n213), .ZN(G45));
  INV_X1    g514(.A(new_n671), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n634), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n664), .A2(new_n666), .A3(new_n657), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  OAI21_X1  g518(.A(new_n190), .B1(new_n269), .B2(new_n278), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  INV_X1    g520(.A(new_n191), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(new_n279), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n605), .A2(new_n635), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND3_X1  g526(.A1(new_n605), .A2(new_n642), .A3(new_n709), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n604), .A2(new_n415), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n708), .A2(new_n608), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n666), .A4(new_n657), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n616), .A2(G472), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n570), .B(new_n578), .C1(new_n595), .C2(new_n551), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n587), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n719), .B1(new_n547), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n723), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(KEYINPUT104), .A3(new_n540), .A4(new_n546), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n708), .A2(new_n620), .A3(new_n676), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NAND4_X1  g544(.A1(new_n716), .A2(new_n665), .A3(new_n702), .A4(new_n725), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  OAI21_X1  g546(.A(new_n264), .B1(new_n285), .B2(KEYINPUT79), .ZN(new_n733));
  INV_X1    g547(.A(new_n265), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n286), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n281), .ZN(new_n736));
  INV_X1    g550(.A(G469), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(KEYINPUT105), .A3(G902), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n288), .B2(KEYINPUT105), .ZN(new_n740));
  INV_X1    g554(.A(new_n279), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n707), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n267), .B1(new_n251), .B2(new_n252), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n270), .B1(new_n745), .B2(new_n265), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n190), .B1(new_n746), .B2(new_n281), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n747), .B2(G469), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n279), .B1(new_n748), .B2(new_n739), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n750), .A3(new_n707), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n484), .A2(new_n418), .A3(new_n487), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n743), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n605), .A3(new_n702), .A4(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n752), .B1(new_n742), .B2(KEYINPUT106), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n605), .A3(new_n702), .A4(new_n751), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n605), .A3(new_n673), .A4(new_n751), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n287), .B2(KEYINPUT45), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n746), .A2(new_n770), .A3(new_n281), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n287), .A2(KEYINPUT45), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n746), .B2(new_n281), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT108), .A4(G469), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(KEYINPUT109), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n772), .A2(new_n775), .B1(G469), .B2(G902), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n741), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n633), .B(new_n361), .C1(new_n621), .C2(new_n622), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n616), .B(new_n617), .Z(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(new_n665), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n785), .A2(new_n707), .A3(new_n682), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT44), .A4(new_n665), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n795), .A3(new_n753), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n795), .B1(new_n794), .B2(new_n753), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n257), .ZN(G39));
  NAND3_X1  g614(.A1(new_n604), .A2(new_n702), .A3(new_n753), .ZN(new_n801));
  INV_X1    g615(.A(new_n547), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n785), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n785), .B2(new_n707), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(new_n407), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n788), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n724), .B2(new_n726), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n753), .ZN(new_n812));
  INV_X1    g626(.A(new_n806), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n804), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n706), .A2(new_n279), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n707), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n812), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n687), .A2(new_n419), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n818), .A2(KEYINPUT117), .A3(new_n708), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT117), .B1(new_n818), .B2(new_n708), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n811), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT50), .Z(new_n822));
  NAND2_X1  g636(.A1(new_n709), .A2(new_n753), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n823), .A2(new_n547), .A3(new_n407), .A4(new_n697), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n623), .A2(new_n633), .ZN(new_n825));
  INV_X1    g639(.A(new_n665), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n723), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n823), .A2(new_n810), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n824), .A2(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n817), .A2(new_n822), .A3(KEYINPUT51), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n634), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(G952), .A3(new_n194), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n605), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT48), .Z(new_n835));
  AOI211_X1 g649(.A(new_n833), .B(new_n835), .C1(new_n716), .C2(new_n811), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n822), .A2(new_n829), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n816), .B1(new_n814), .B2(KEYINPUT116), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(KEYINPUT116), .B2(new_n814), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n839), .B2(new_n812), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n830), .B(new_n836), .C1(new_n840), .C2(KEYINPUT51), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n749), .A2(new_n540), .A3(new_n707), .A4(new_n651), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n697), .A2(new_n677), .A3(new_n488), .A4(new_n671), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n586), .A2(KEYINPUT32), .A3(new_n587), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT32), .B1(new_n586), .B2(new_n587), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(new_n695), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n685), .A2(new_n418), .A3(new_n623), .A4(new_n639), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n848), .A2(new_n849), .A3(new_n701), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  INV_X1    g665(.A(new_n739), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n735), .A2(new_n736), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n737), .B1(new_n853), .B2(new_n190), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n854), .B2(new_n744), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n191), .B1(new_n855), .B2(new_n279), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n851), .A3(new_n856), .A4(new_n826), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n845), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n674), .A2(new_n703), .A3(new_n731), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n842), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n857), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n603), .A2(new_n673), .A3(new_n488), .A4(new_n289), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n603), .A2(new_n702), .A3(new_n488), .A4(new_n289), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n660), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT52), .A4(new_n731), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n860), .A2(KEYINPUT113), .A3(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT111), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n358), .A2(new_n361), .A3(new_n639), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n490), .A2(new_n869), .A3(new_n411), .A4(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n609), .A2(new_n610), .A3(new_n871), .A4(new_n411), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT111), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n619), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n619), .A2(new_n490), .A3(new_n411), .A4(new_n831), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n661), .A2(new_n613), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n605), .B(new_n709), .C1(new_n635), .C2(new_n642), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n729), .A2(new_n717), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n289), .A2(new_n603), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n641), .A2(new_n405), .A3(new_n413), .A4(new_n671), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n752), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n660), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n665), .A2(new_n725), .A3(new_n702), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n759), .A2(new_n885), .A3(new_n751), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n766), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n763), .B2(new_n758), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n880), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n860), .A2(new_n865), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n880), .A3(new_n888), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n868), .A2(new_n890), .B1(KEYINPUT53), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n889), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n878), .A2(new_n717), .ZN(new_n897));
  INV_X1    g711(.A(new_n728), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n724), .B2(new_n726), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n729), .A2(KEYINPUT114), .A3(new_n717), .A4(new_n878), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n877), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n766), .A2(new_n884), .A3(new_n886), .A4(KEYINPUT53), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n763), .B2(new_n758), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n866), .A3(new_n867), .A4(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  OAI22_X1  g722(.A1(new_n841), .A2(new_n908), .B1(G952), .B2(G953), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n688), .A2(new_n419), .A3(new_n191), .A4(new_n786), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n697), .B1(new_n815), .B2(KEYINPUT49), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n802), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n194), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n190), .B1(new_n895), .B2(new_n905), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n448), .A2(new_n459), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n457), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n895), .A2(new_n905), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n925), .A3(G210), .A4(G902), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n921), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n917), .B2(G210), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n924), .A2(G210), .A3(G902), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT118), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(KEYINPUT119), .A3(new_n926), .A4(new_n928), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n922), .B1(new_n931), .B2(new_n934), .ZN(G51));
  INV_X1    g749(.A(new_n907), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n906), .B1(new_n895), .B2(new_n905), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n777), .B(KEYINPUT57), .ZN(new_n939));
  OAI22_X1  g753(.A1(new_n938), .A2(new_n939), .B1(new_n269), .B2(new_n278), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n917), .A2(new_n772), .A3(new_n775), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n915), .B1(new_n940), .B2(new_n941), .ZN(G54));
  NAND2_X1  g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT120), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n190), .B(new_n945), .C1(new_n895), .C2(new_n905), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n916), .B1(new_n946), .B2(new_n354), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n924), .A2(G902), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n948), .A2(new_n356), .A3(new_n945), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT121), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n356), .B1(new_n948), .B2(new_n945), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n354), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n916), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(G60));
  INV_X1    g769(.A(new_n631), .ZN(new_n956));
  XNOR2_X1  g770(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n916), .B1(new_n938), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n908), .B2(new_n959), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n895), .B2(new_n905), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n916), .B1(new_n966), .B2(new_n544), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n648), .B(new_n965), .C1(new_n895), .C2(new_n905), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n408), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n880), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n919), .B1(G898), .B2(new_n194), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  XNOR2_X1  g791(.A(new_n568), .B(new_n343), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n752), .B1(new_n870), .B2(new_n634), .ZN(new_n979));
  AND4_X1   g793(.A1(new_n605), .A2(new_n289), .A3(new_n682), .A4(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n793), .ZN(new_n981));
  INV_X1    g795(.A(new_n798), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n674), .A2(new_n703), .A3(new_n731), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n984), .B(KEYINPUT62), .C1(new_n698), .C2(new_n681), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n699), .B2(new_n859), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n983), .A2(new_n988), .A3(new_n807), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n978), .B1(new_n989), .B2(G953), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n984), .B1(new_n793), .B2(new_n798), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(KEYINPUT123), .B(new_n984), .C1(new_n793), .C2(new_n798), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n803), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n813), .B2(new_n804), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n547), .A2(new_n604), .A3(new_n849), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n785), .A2(new_n707), .A3(new_n682), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n764), .A2(new_n766), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n667), .B1(new_n1002), .B2(new_n194), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n990), .B1(new_n1003), .B2(new_n978), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT124), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G72));
  NAND3_X1  g821(.A1(new_n995), .A2(new_n1001), .A3(new_n880), .ZN(new_n1008));
  XNOR2_X1  g822(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n600), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n584), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1014), .A2(new_n692), .A3(new_n1011), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n915), .B1(new_n893), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n983), .A2(new_n988), .A3(new_n807), .A4(new_n880), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n1011), .ZN(new_n1022));
  INV_X1    g836(.A(new_n692), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g838(.A(KEYINPUT126), .B(new_n692), .C1(new_n1021), .C2(new_n1011), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT127), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n890), .A2(new_n867), .A3(new_n866), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n892), .A2(KEYINPUT53), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1028), .A2(new_n1029), .A3(new_n1017), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n916), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1014), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n692), .B1(new_n1021), .B2(new_n1011), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(new_n1020), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT127), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1027), .A2(new_n1037), .ZN(G57));
endmodule


