//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(KEYINPUT66), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n190), .A2(new_n192), .B1(KEYINPUT2), .B2(G113), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n193), .A2(KEYINPUT67), .A3(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n193), .A2(new_n198), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT30), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G137), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n207), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(new_n208), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT64), .A3(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  AND4_X1   g042(.A1(KEYINPUT65), .A2(new_n225), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n223), .A2(G146), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n222), .B2(new_n224), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT65), .B1(new_n231), .B2(new_n228), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n223), .B2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(G146), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n234), .A2(G128), .B1(new_n226), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n219), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT0), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n227), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n226), .A2(new_n235), .B1(KEYINPUT0), .B2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n227), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n239), .A2(new_n231), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n213), .A2(new_n208), .A3(new_n215), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n217), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n206), .B1(new_n237), .B2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n223), .A2(KEYINPUT64), .A3(G146), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT64), .B1(new_n223), .B2(G146), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n226), .B(new_n228), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n236), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n246), .B(new_n206), .C1(new_n254), .C2(new_n218), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n205), .B1(new_n247), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n193), .A2(new_n198), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n201), .B2(new_n202), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(new_n246), .C1(new_n254), .C2(new_n218), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(G101), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n262), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n246), .B1(new_n254), .B2(new_n218), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n205), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n237), .A2(KEYINPUT28), .A3(new_n259), .A4(new_n246), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n265), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n257), .A2(new_n276), .A3(new_n260), .A4(new_n265), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n278), .A2(KEYINPUT68), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT68), .B1(new_n278), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n187), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n187), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n260), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n274), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n269), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(KEYINPUT70), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n270), .A2(KEYINPUT30), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n259), .B1(new_n298), .B2(new_n255), .ZN(new_n299));
  INV_X1    g113(.A(new_n260), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n274), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(new_n290), .C1(new_n274), .C2(new_n273), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(G472), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n304), .B1(new_n303), .B2(G472), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n282), .B(new_n285), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT9), .B(G234), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n309), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G104), .B(G107), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT80), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G104), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G107), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G101), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(new_n315), .B2(G107), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n317), .A3(G104), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n322), .A2(new_n324), .A3(new_n313), .A4(new_n316), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n314), .B(new_n321), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n254), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n322), .A2(new_n324), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(KEYINPUT78), .A3(new_n313), .A4(new_n316), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n326), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n324), .A3(new_n316), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G101), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n334), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(G101), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n330), .A2(KEYINPUT10), .B1(new_n341), .B2(new_n242), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  INV_X1    g157(.A(new_n231), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n234), .A2(KEYINPUT81), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n226), .A2(new_n346), .A3(KEYINPUT1), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(G128), .A3(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n252), .A2(new_n253), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n329), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n245), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT82), .B(new_n343), .C1(new_n329), .C2(new_n349), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n342), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n329), .A2(new_n254), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n314), .A2(new_n321), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n333), .B2(new_n332), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n344), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n229), .B2(new_n232), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n353), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(KEYINPUT12), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(KEYINPUT12), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n355), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G110), .B(G140), .ZN(new_n366));
  INV_X1    g180(.A(G953), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(G227), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n366), .B(new_n368), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n341), .A2(new_n242), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n330), .A2(KEYINPUT10), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n352), .A2(new_n372), .A3(new_n373), .A4(new_n354), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT83), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n342), .A2(new_n352), .A3(new_n376), .A4(new_n354), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n353), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n355), .A2(new_n369), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n371), .B(G469), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n355), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n370), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n363), .A2(new_n364), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n379), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n293), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n311), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n194), .A2(KEYINPUT72), .A3(G128), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT72), .B1(new_n194), .B2(G128), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n393), .A2(new_n394), .B1(new_n194), .B2(G128), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT24), .B(G110), .Z(new_n396));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(G119), .B2(new_n227), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n194), .A2(KEYINPUT23), .A3(G128), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n398), .A2(new_n399), .B1(G119), .B2(new_n227), .ZN(new_n400));
  OAI22_X1  g214(.A1(new_n395), .A2(new_n396), .B1(new_n400), .B2(G110), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT73), .A2(G125), .ZN(new_n402));
  NOR2_X1   g216(.A1(KEYINPUT73), .A2(G125), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G125), .A2(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n404), .B2(G140), .ZN(new_n409));
  OAI211_X1 g223(.A(G146), .B(new_n407), .C1(new_n409), .C2(new_n405), .ZN(new_n410));
  XOR2_X1   g224(.A(G125), .B(G140), .Z(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(G146), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(KEYINPUT73), .A2(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT73), .A2(G125), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(G140), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n408), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n405), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR4_X1   g232(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT16), .A4(G140), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n221), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n410), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n395), .A2(new_n396), .B1(new_n400), .B2(G110), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT74), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n413), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n367), .A2(G221), .A3(G234), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT22), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n214), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT75), .Z(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(new_n413), .C1(new_n423), .C2(new_n424), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT76), .B1(new_n432), .B2(KEYINPUT25), .ZN(new_n433));
  INV_X1    g247(.A(new_n413), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n416), .A2(new_n417), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT16), .ZN(new_n436));
  AOI21_X1  g250(.A(G146), .B1(new_n436), .B2(new_n407), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n418), .A2(new_n221), .A3(new_n419), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n422), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n422), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n434), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n428), .B(KEYINPUT75), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n431), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT25), .A3(new_n293), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT77), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n293), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT76), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n432), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n433), .A2(new_n448), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G217), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G234), .B2(new_n293), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G902), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n454), .A2(new_n456), .B1(new_n445), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n263), .A2(G214), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(G143), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n223), .A2(KEYINPUT88), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(G214), .A4(new_n263), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT17), .A4(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n420), .A2(new_n410), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT90), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n461), .A2(new_n464), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(G131), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n420), .A2(new_n410), .A3(new_n472), .A4(new_n465), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n412), .B1(new_n435), .B2(new_n221), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n476), .A2(new_n468), .A3(KEYINPUT18), .A4(G131), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n468), .A2(new_n476), .B1(KEYINPUT18), .B2(G131), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n315), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(new_n482), .A3(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n293), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G475), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n409), .A2(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(KEYINPUT19), .B2(new_n411), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n410), .B1(new_n493), .B2(G146), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n479), .B1(new_n494), .B2(new_n469), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n483), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n491), .B1(new_n485), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT20), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n485), .A2(new_n496), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT20), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n490), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n489), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n309), .A2(new_n455), .A3(G953), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT13), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n227), .B2(G143), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n223), .A2(G128), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT92), .A3(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n227), .A2(G143), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n223), .A2(KEYINPUT13), .A3(G128), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G134), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n514), .A3(new_n207), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n196), .A2(G122), .ZN(new_n519));
  INV_X1    g333(.A(G122), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G116), .ZN(new_n521));
  OR3_X1    g335(.A1(new_n519), .A2(new_n521), .A3(G107), .ZN(new_n522));
  OAI21_X1  g336(.A(G107), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT93), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n517), .A2(new_n524), .A3(new_n527), .A4(new_n518), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n512), .A2(new_n514), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G134), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n518), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(new_n520), .B2(G116), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT94), .ZN(new_n535));
  INV_X1    g349(.A(new_n519), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(KEYINPUT14), .C1(new_n520), .C2(G116), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g355(.A1(new_n520), .A2(KEYINPUT14), .A3(G116), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(KEYINPUT95), .A3(new_n536), .A4(new_n538), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n533), .B1(new_n544), .B2(G107), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n507), .B1(new_n529), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(G107), .ZN(new_n547));
  INV_X1    g361(.A(new_n533), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(new_n526), .A3(new_n528), .A4(new_n506), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(KEYINPUT96), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(new_n507), .C1(new_n529), .C2(new_n545), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n293), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(KEYINPUT15), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n554), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n505), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G210), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n205), .A2(new_n341), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT5), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n196), .A2(KEYINPUT5), .A3(G119), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(G113), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT84), .A4(G113), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n201), .A2(new_n202), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n358), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(G110), .B(G122), .Z(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n572), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n205), .A2(new_n341), .B1(new_n569), .B2(new_n358), .ZN(new_n574));
  INV_X1    g388(.A(new_n572), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n242), .A2(new_n404), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n254), .B2(new_n404), .ZN(new_n582));
  INV_X1    g396(.A(G224), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G953), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT86), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n582), .B(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n567), .A2(new_n568), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n203), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT87), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n329), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT87), .B1(new_n569), .B2(new_n358), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n358), .A2(new_n203), .A3(new_n565), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n572), .B(KEYINPUT8), .Z(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n584), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n574), .A2(new_n575), .B1(new_n582), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n596), .B(new_n599), .C1(new_n582), .C2(new_n598), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n293), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n561), .B1(new_n587), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n580), .A2(new_n586), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(new_n293), .A3(new_n560), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G214), .B1(G237), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(G952), .A3(new_n367), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT21), .B(G898), .Z(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n605), .A2(new_n606), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n559), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n307), .A2(new_n392), .A3(new_n458), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AOI21_X1  g433(.A(KEYINPUT82), .B1(new_n361), .B2(new_n343), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n351), .B(KEYINPUT10), .C1(new_n358), .C2(new_n360), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n376), .B1(new_n622), .B2(new_n342), .ZN(new_n623));
  AND4_X1   g437(.A1(new_n376), .A2(new_n342), .A3(new_n352), .A4(new_n354), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n245), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n369), .B1(new_n625), .B2(new_n355), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n388), .B(new_n293), .C1(new_n626), .C2(new_n385), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n391), .A3(new_n380), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n278), .B2(new_n293), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT68), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n283), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n278), .A2(KEYINPUT68), .A3(new_n279), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n458), .A2(new_n628), .A3(new_n310), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT97), .Z(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n551), .A2(new_n637), .A3(new_n553), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n546), .A2(KEYINPUT33), .A3(new_n550), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n293), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G478), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n554), .A2(G478), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n644));
  INV_X1    g458(.A(new_n490), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n502), .A2(KEYINPUT91), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n497), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n504), .B1(new_n647), .B2(new_n503), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n488), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n641), .A2(new_n650), .A3(new_n642), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n644), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n602), .A2(new_n653), .A3(new_n604), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT98), .B(new_n561), .C1(new_n587), .C2(new_n601), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n606), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n652), .A2(new_n656), .A3(new_n614), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n315), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n500), .B2(KEYINPUT20), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n501), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n500), .A2(new_n662), .A3(KEYINPUT20), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n489), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n558), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n614), .A3(new_n656), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n636), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NOR2_X1   g486(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n425), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n457), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n454), .B2(new_n456), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n392), .A2(new_n617), .A3(new_n634), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT37), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G110), .ZN(G12));
  NAND2_X1  g494(.A1(new_n303), .A2(G472), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT71), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n303), .A2(new_n304), .A3(G472), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n632), .A2(new_n633), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n284), .B1(new_n685), .B2(new_n187), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n676), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n628), .A2(new_n310), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n656), .ZN(new_n689));
  OR3_X1    g503(.A1(new_n612), .A2(KEYINPUT102), .A3(G900), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT102), .B1(new_n612), .B2(G900), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n608), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n666), .A2(new_n667), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n687), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XOR2_X1   g510(.A(new_n692), .B(KEYINPUT39), .Z(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n392), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT40), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n605), .B(KEYINPUT38), .Z(new_n701));
  INV_X1    g515(.A(new_n606), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n287), .A2(new_n288), .A3(new_n274), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n266), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n293), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n266), .B2(new_n706), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n282), .A2(new_n285), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n558), .B1(new_n648), .B2(new_n488), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n676), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n703), .A2(new_n704), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n704), .B1(new_n703), .B2(new_n714), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n700), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT105), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n223), .ZN(G45));
  INV_X1    g533(.A(new_n692), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n652), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n687), .A2(new_n689), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  INV_X1    g537(.A(new_n458), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n684), .B2(new_n686), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n383), .A2(new_n386), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n293), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n728), .A2(new_n310), .A3(new_n627), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(new_n657), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND3_X1  g546(.A1(new_n669), .A2(new_n725), .A3(new_n729), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NAND3_X1  g548(.A1(new_n728), .A2(new_n310), .A3(new_n627), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n656), .ZN(new_n736));
  INV_X1    g550(.A(new_n559), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n687), .A2(new_n736), .A3(new_n737), .A4(new_n615), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  INV_X1    g553(.A(new_n630), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n267), .A2(new_n277), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n265), .B1(new_n289), .B2(new_n269), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n279), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n724), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n736), .A2(new_n615), .A3(new_n712), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT106), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR2_X1   g562(.A1(new_n744), .A2(new_n676), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n736), .A2(new_n721), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NOR2_X1   g565(.A1(new_n605), .A2(new_n702), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n628), .A2(new_n310), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n307), .A3(new_n458), .A4(new_n721), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n641), .A2(new_n650), .A3(new_n642), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n650), .B1(new_n641), .B2(new_n642), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n752), .A3(new_n649), .A4(new_n692), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n688), .A3(new_n755), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n284), .B1(new_n682), .B2(new_n683), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n283), .A2(new_n187), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n724), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n754), .A2(new_n755), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n216), .ZN(G33));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n693), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n666), .A2(KEYINPUT107), .A3(new_n667), .A4(new_n692), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n725), .A2(new_n767), .A3(new_n753), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  OAI21_X1  g584(.A(new_n371), .B1(new_n378), .B2(new_n379), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT108), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n773), .A2(new_n777), .A3(G469), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n391), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n391), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n785), .A3(KEYINPUT46), .A4(new_n391), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n781), .A2(new_n784), .A3(new_n627), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n310), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n697), .ZN(new_n789));
  INV_X1    g603(.A(new_n752), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n758), .A2(new_n505), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n758), .A2(KEYINPUT43), .A3(new_n505), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n634), .B(new_n676), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n791), .B1(new_n796), .B2(KEYINPUT44), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  INV_X1    g612(.A(new_n634), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n677), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(KEYINPUT110), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n796), .A2(KEYINPUT44), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n789), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT111), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n214), .ZN(G39));
  NOR3_X1   g621(.A1(new_n307), .A2(new_n759), .A3(new_n458), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n310), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT47), .B1(new_n787), .B2(new_n310), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NOR3_X1   g626(.A1(new_n735), .A2(new_n608), .A3(new_n790), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n686), .A2(new_n813), .A3(new_n458), .A4(new_n710), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n649), .A3(new_n758), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n798), .A2(new_n609), .A3(new_n745), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n736), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n817), .A3(G952), .A4(new_n367), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT117), .Z(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n788), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n787), .A2(KEYINPUT47), .A3(new_n310), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n728), .A2(new_n627), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n310), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n752), .B(new_n816), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n798), .A2(new_n609), .A3(new_n729), .A4(new_n745), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n701), .A2(new_n702), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT50), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n798), .A2(new_n813), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT116), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n749), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n814), .B(new_n505), .C1(new_n757), .C2(new_n756), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n819), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  INV_X1    g655(.A(new_n656), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n392), .A2(new_n842), .A3(new_n711), .A4(new_n713), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT113), .B1(new_n843), .B2(new_n720), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n714), .A2(new_n689), .A3(new_n845), .A4(new_n692), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n695), .A2(new_n722), .A3(new_n750), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT52), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n649), .B1(new_n756), .B2(new_n757), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(KEYINPUT112), .A3(new_n559), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n652), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n616), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n635), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n618), .A3(new_n678), .ZN(new_n857));
  INV_X1    g671(.A(new_n769), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n764), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n733), .A2(new_n738), .A3(new_n730), .A4(new_n746), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n667), .A2(new_n720), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n307), .A2(new_n666), .A3(new_n677), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n721), .A2(new_n749), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n753), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n695), .A2(new_n722), .A3(new_n750), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n844), .A2(new_n846), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n849), .A2(new_n859), .A3(new_n866), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n856), .A2(new_n618), .A3(new_n678), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n754), .A2(new_n755), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n760), .A2(new_n763), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n877), .A3(new_n769), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n746), .A2(new_n730), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n729), .A2(new_n307), .A3(new_n458), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n735), .A2(new_n559), .A3(new_n614), .A4(new_n656), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n880), .A2(new_n669), .B1(new_n881), .B2(new_n687), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n864), .A2(new_n753), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n870), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n841), .B1(new_n873), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT114), .B1(new_n871), .B2(new_n872), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n873), .A2(new_n890), .A3(new_n886), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT115), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n873), .A2(new_n886), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n832), .A2(new_n763), .ZN(new_n896));
  NOR2_X1   g710(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n897));
  AND2_X1   g711(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n840), .A2(new_n889), .A3(new_n895), .A4(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n824), .B(KEYINPUT49), .Z(new_n903));
  NOR4_X1   g717(.A1(new_n792), .A2(new_n711), .A3(new_n702), .A4(new_n311), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n458), .A3(new_n701), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n367), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n293), .B1(new_n873), .B2(new_n886), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n909), .B2(G210), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n580), .A2(new_n586), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n587), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n873), .A2(new_n886), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(G902), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT119), .B(new_n293), .C1(new_n873), .C2(new_n886), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n561), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n914), .B1(new_n920), .B2(new_n922), .ZN(G51));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n924));
  INV_X1    g738(.A(new_n779), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n390), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n873), .A2(new_n890), .A3(new_n886), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n890), .B1(new_n873), .B2(new_n886), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n919), .A2(new_n925), .B1(new_n930), .B2(new_n726), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n924), .B1(new_n931), .B2(new_n907), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n930), .A2(new_n726), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n917), .A2(new_n918), .A3(new_n779), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT121), .B(new_n908), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(G54));
  NAND3_X1  g750(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n498), .A2(new_n499), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n938), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .A4(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n939), .A2(new_n908), .A3(new_n941), .ZN(G60));
  INV_X1    g756(.A(new_n929), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n891), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n638), .A2(new_n639), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n555), .A2(new_n293), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n944), .A2(new_n952), .A3(new_n945), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n948), .B1(new_n895), .B2(new_n889), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n908), .B1(new_n955), .B2(new_n945), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n916), .A2(new_n674), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n916), .A2(new_n959), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n908), .B(new_n960), .C1(new_n961), .C2(new_n445), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n611), .B2(new_n583), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n860), .A2(new_n857), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  INV_X1    g780(.A(new_n580), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(G898), .B2(new_n367), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  INV_X1    g783(.A(new_n717), .ZN(new_n970));
  NAND2_X1  g784(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n867), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n717), .B2(new_n848), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n805), .A2(new_n811), .A3(new_n972), .A4(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n725), .A2(new_n854), .A3(new_n698), .A4(new_n753), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n367), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n247), .A2(new_n256), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n493), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g798(.A1(G900), .A2(G953), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n805), .A2(new_n811), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n763), .A2(new_n712), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n787), .A2(new_n310), .A3(new_n698), .A4(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n877), .B(new_n867), .C1(new_n988), .C2(new_n656), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n769), .A3(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n981), .B(new_n985), .C1(new_n991), .C2(G953), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n979), .A2(new_n993), .A3(new_n982), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n984), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n367), .B1(G227), .B2(G900), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n996), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n984), .A2(new_n998), .A3(new_n992), .A4(new_n994), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G72));
  NOR2_X1   g814(.A1(new_n299), .A2(new_n300), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(new_n274), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n965), .ZN(new_n1004));
  OR3_X1    g818(.A1(new_n976), .A2(new_n1004), .A3(new_n978), .ZN(new_n1005));
  XNOR2_X1  g819(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n629), .A2(new_n293), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n1003), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n887), .A2(new_n888), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1008), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1010), .A2(new_n1011), .A3(new_n1002), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1001), .A2(new_n274), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n986), .A2(new_n769), .A3(new_n965), .A4(new_n990), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1013), .B1(new_n1015), .B2(new_n1008), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1014), .B1(new_n1016), .B2(new_n907), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1013), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n805), .A2(new_n811), .A3(new_n769), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1019), .A2(new_n1004), .A3(new_n989), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1018), .B1(new_n1020), .B2(new_n1011), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(KEYINPUT127), .A3(new_n908), .ZN(new_n1022));
  AOI221_X4 g836(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .C1(new_n1017), .C2(new_n1022), .ZN(G57));
endmodule


