//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XNOR2_X1  g0005(.A(KEYINPUT65), .B(G238), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(new_n207), .A2(G68), .B1(G77), .B2(G244), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G58), .A2(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AND2_X1   g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n202), .A2(new_n217), .ZN(new_n218));
  NOR4_X1   g0018(.A1(new_n212), .A2(new_n213), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G87), .A2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n219), .A2(new_n220), .B1(G1), .B2(G20), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT64), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n226), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT66), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n224), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n249), .A2(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n227), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(KEYINPUT67), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n225), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n258), .A2(new_n263), .B1(new_n202), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G50), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G222), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n276), .C1(G77), .C2(new_n271), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n276), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n278), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n277), .B(new_n281), .C1(new_n217), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n284), .A2(G179), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n270), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n271), .A2(G232), .A3(new_n273), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G107), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(new_n292), .A3(G1698), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n206), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n276), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n283), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G244), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n300), .A3(new_n281), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n289), .B(new_n294), .C1(new_n206), .C2(new_n296), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n280), .B1(new_n304), .B2(new_n276), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT69), .B1(new_n305), .B2(new_n300), .ZN(new_n306));
  OAI21_X1  g0106(.A(G190), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n302), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(KEYINPUT69), .A3(new_n300), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G200), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n252), .B(KEYINPUT70), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n311), .A2(new_n249), .B1(new_n250), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n224), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n263), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n266), .A2(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n268), .A2(G77), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n307), .A2(new_n310), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT9), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n270), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n284), .A2(G200), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n267), .A2(KEYINPUT9), .A3(new_n269), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n284), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT10), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n288), .B(new_n322), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n290), .A2(new_n292), .A3(G226), .A4(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT76), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n271), .A2(new_n335), .A3(G226), .A4(G1698), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n290), .A2(new_n292), .A3(G223), .A4(new_n273), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G87), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT77), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n340), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n334), .A4(new_n336), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n276), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n280), .B1(new_n299), .B2(G232), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n285), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT78), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n345), .A2(new_n352), .A3(new_n346), .A4(new_n347), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n291), .A2(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT73), .ZN(new_n361));
  AOI21_X1  g0161(.A(G20), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT74), .B1(new_n362), .B2(KEYINPUT7), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT73), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT73), .B1(new_n290), .B2(new_n292), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n224), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G68), .ZN(new_n372));
  XNOR2_X1  g0172(.A(G58), .B(G68), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(KEYINPUT16), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT75), .B1(new_n291), .B2(G33), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n380), .A3(new_n292), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n369), .B1(new_n271), .B2(G20), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n374), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n376), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n375), .A2(new_n263), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n249), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n266), .ZN(new_n389));
  INV_X1    g0189(.A(new_n268), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n388), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT79), .A4(new_n353), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n356), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n356), .A2(new_n393), .A3(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n332), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n345), .A2(G190), .A3(new_n347), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n350), .A2(G200), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n387), .A2(new_n392), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n263), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n385), .B1(new_n371), .B2(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n391), .B1(new_n408), .B2(new_n386), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n401), .A4(new_n402), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n308), .A2(new_n309), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n320), .B1(new_n412), .B2(new_n346), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n308), .A2(new_n285), .A3(new_n309), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n290), .A2(new_n292), .A3(G232), .A4(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT71), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n271), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n271), .A2(G226), .A3(new_n273), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n280), .B1(new_n422), .B2(new_n276), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n299), .A2(G238), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  OAI21_X1  g0227(.A(G169), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT14), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G179), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(G169), .C1(new_n426), .C2(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n268), .A2(G68), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT72), .Z(new_n436));
  OAI22_X1  g0236(.A1(new_n253), .A2(new_n202), .B1(new_n224), .B2(G68), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n250), .A2(new_n314), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n263), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT11), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n266), .A2(new_n377), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n415), .B1(new_n434), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n430), .A2(G190), .ZN(new_n447));
  INV_X1    g0247(.A(G200), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n444), .C1(new_n448), .C2(new_n430), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n411), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n400), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n224), .C1(G33), .C2(new_n214), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n263), .B(new_n453), .C1(new_n224), .C2(G116), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n266), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n265), .B1(G1), .B2(new_n260), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n263), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G116), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT84), .ZN(new_n463));
  INV_X1    g0263(.A(G41), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(KEYINPUT84), .B2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n282), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G270), .ZN(new_n473));
  INV_X1    g0273(.A(G303), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n296), .A2(new_n211), .B1(new_n271), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n293), .A2(new_n215), .A3(G1698), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n276), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(G274), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n462), .B1(G200), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n479), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G190), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n210), .A2(G20), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT23), .ZN(new_n486));
  INV_X1    g0286(.A(new_n250), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(G116), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n271), .A2(new_n224), .A3(G87), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT90), .B(KEYINPUT22), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT24), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n263), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n460), .A2(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT91), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT25), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n265), .C2(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n265), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(KEYINPUT91), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT92), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT92), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n498), .A2(new_n507), .A3(new_n501), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n497), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n472), .A2(G264), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n290), .A2(new_n292), .A3(G250), .A4(new_n273), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n296), .C2(new_n215), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n276), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n511), .A2(new_n515), .A3(new_n478), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n285), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n346), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n462), .A2(G169), .A3(new_n479), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n462), .A2(G179), .A3(new_n481), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n462), .A2(KEYINPUT21), .A3(G169), .A4(new_n479), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n460), .A2(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n266), .A2(new_n214), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n210), .B1(new_n382), .B2(new_n383), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n253), .A2(new_n314), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n214), .A2(new_n210), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n224), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n530), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n528), .B(new_n529), .C1(new_n538), .C2(new_n406), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n290), .A2(new_n292), .A3(G244), .A4(new_n273), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n271), .A2(KEYINPUT81), .A3(G244), .A4(new_n273), .ZN(new_n543));
  XOR2_X1   g0343(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n452), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n290), .A2(new_n292), .A3(new_n273), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT4), .A4(G244), .ZN(new_n549));
  INV_X1    g0349(.A(new_n296), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G250), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT83), .B1(new_n540), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n276), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n478), .B1(new_n471), .B2(new_n215), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT85), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT85), .B(new_n478), .C1(new_n471), .C2(new_n215), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n560), .A3(new_n346), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n540), .A2(new_n552), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n548), .B1(new_n550), .B2(G250), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n452), .A3(new_n553), .A4(new_n545), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n556), .B1(new_n564), .B2(new_n276), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n539), .B(new_n561), .C1(G169), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT86), .ZN(new_n567));
  INV_X1    g0367(.A(new_n556), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n555), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n285), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n561), .A4(new_n539), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n517), .A2(G200), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n516), .A2(G190), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n509), .A3(new_n497), .A4(new_n575), .ZN(new_n576));
  OR2_X1    g0376(.A1(G238), .A2(G1698), .ZN(new_n577));
  INV_X1    g0377(.A(G244), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n290), .A2(new_n577), .A3(new_n292), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G116), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n581), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n276), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n469), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n282), .A2(G250), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n469), .A2(G274), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n312), .A2(new_n266), .ZN(new_n593));
  INV_X1    g0393(.A(G87), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n263), .A2(new_n459), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n487), .A2(new_n596), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n534), .A2(new_n594), .B1(new_n421), .B2(new_n224), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n596), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n271), .A2(new_n224), .A3(G68), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT88), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n271), .A2(new_n602), .A3(new_n224), .A4(G68), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n593), .B(new_n595), .C1(new_n604), .C2(new_n263), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n592), .B(new_n605), .C1(new_n327), .C2(new_n591), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n593), .B1(new_n604), .B2(new_n263), .ZN(new_n607));
  XOR2_X1   g0407(.A(new_n312), .B(KEYINPUT89), .Z(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n460), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n591), .A2(new_n285), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n586), .A2(new_n346), .A3(new_n590), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n606), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n569), .A2(new_n327), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n448), .B1(new_n555), .B2(new_n560), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n616), .A2(new_n539), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n573), .A2(new_n576), .A3(new_n615), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n451), .A2(new_n484), .A3(new_n527), .A4(new_n621), .ZN(G372));
  INV_X1    g0422(.A(KEYINPUT93), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n330), .A2(new_n331), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n434), .A2(new_n445), .ZN(new_n626));
  INV_X1    g0426(.A(new_n415), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n405), .A3(new_n410), .A4(new_n449), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT18), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n409), .B2(new_n354), .ZN(new_n631));
  INV_X1    g0431(.A(new_n354), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n393), .A2(new_n632), .A3(KEYINPUT18), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n625), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n623), .B1(new_n635), .B2(new_n288), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n405), .A2(new_n410), .A3(new_n449), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n446), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n624), .ZN(new_n639));
  INV_X1    g0439(.A(new_n288), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(KEYINPUT93), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n618), .B1(new_n567), .B2(new_n572), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(new_n526), .A3(new_n576), .A4(new_n615), .ZN(new_n644));
  INV_X1    g0444(.A(new_n566), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n615), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n614), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n567), .A2(new_n615), .A3(new_n572), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n644), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n451), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(G369));
  INV_X1    g0453(.A(G13), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n264), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n520), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n510), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n576), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n520), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n462), .A2(new_n661), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n667), .B(new_n668), .Z(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n484), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n661), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(new_n662), .ZN(G399));
  INV_X1    g0475(.A(new_n228), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n534), .A2(new_n594), .A3(new_n457), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n223), .B2(new_n678), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT97), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n567), .A2(new_n646), .A3(new_n615), .A4(new_n572), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n606), .A2(new_n614), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n687), .B2(new_n566), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n614), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n686), .A2(KEYINPUT96), .A3(new_n614), .A4(new_n688), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n644), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n685), .B1(new_n693), .B2(new_n672), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n651), .A2(new_n685), .A3(new_n672), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n586), .A2(new_n515), .A3(new_n511), .A4(new_n590), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n473), .A2(new_n477), .A3(G179), .A4(new_n478), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n555), .B(new_n568), .C1(new_n699), .C2(KEYINPUT30), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n516), .B1(new_n555), .B2(new_n560), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n346), .A3(new_n479), .A4(new_n591), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n701), .A2(new_n702), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n699), .A3(new_n565), .A4(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT31), .B1(new_n710), .B2(new_n661), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(KEYINPUT95), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n661), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n712), .B1(new_n717), .B2(KEYINPUT95), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n621), .A2(new_n484), .A3(new_n527), .A4(new_n672), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n698), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n684), .B1(new_n697), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n697), .A2(new_n684), .A3(new_n721), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n683), .B1(new_n725), .B2(G1), .ZN(G364));
  INV_X1    g0526(.A(new_n670), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n698), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n655), .A2(G45), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n678), .A2(G1), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n671), .A3(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n225), .B1(G20), .B2(new_n285), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n224), .A2(new_n346), .A3(new_n327), .A4(G200), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT100), .ZN(new_n737));
  INV_X1    g0537(.A(G58), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n271), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n346), .A2(G200), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT101), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G190), .A2(G200), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G20), .A3(new_n346), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT32), .B1(new_n747), .B2(G159), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n747), .A2(KEYINPUT32), .A3(G159), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n744), .A2(new_n210), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n224), .A2(new_n346), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n739), .B(new_n750), .C1(G68), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n327), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n224), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G97), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n752), .A2(new_n327), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G50), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n742), .A2(new_n327), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n745), .A2(G20), .A3(G179), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n761), .A2(G87), .B1(G77), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n754), .A2(new_n758), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT102), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n761), .A2(G303), .B1(G311), .B2(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  INV_X1    g0568(.A(new_n736), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n747), .A2(G329), .ZN(new_n771));
  XOR2_X1   g0571(.A(KEYINPUT33), .B(G317), .Z(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT103), .ZN(new_n773));
  INV_X1    g0573(.A(new_n753), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n770), .A2(new_n271), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n759), .A2(G326), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n756), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G283), .B2(new_n743), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n735), .B1(new_n766), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n735), .A2(new_n733), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n223), .A2(G45), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n365), .A2(new_n366), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n228), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(G45), .C2(new_n243), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n271), .A2(new_n228), .ZN(new_n788));
  INV_X1    g0588(.A(G355), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n788), .A2(new_n789), .B1(G116), .B2(new_n228), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n782), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n734), .A2(new_n781), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n732), .A2(new_n793), .ZN(G396));
  NAND2_X1  g0594(.A1(new_n651), .A2(new_n672), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n319), .A2(new_n661), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n321), .A2(new_n796), .B1(new_n413), .B2(new_n414), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n413), .A2(new_n414), .A3(new_n672), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT105), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT105), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n319), .B1(new_n412), .B2(G190), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(new_n310), .B1(new_n319), .B2(new_n661), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n798), .C1(new_n803), .C2(new_n415), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n800), .A2(new_n804), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n651), .A2(new_n807), .A3(new_n672), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(new_n720), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n731), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n731), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n759), .A2(G303), .B1(G311), .B2(new_n747), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n774), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n744), .A2(new_n594), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n761), .A2(G107), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n271), .B1(new_n763), .B2(G116), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n758), .A4(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n817), .B(new_n822), .C1(G294), .C2(new_n736), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n785), .B1(new_n761), .B2(G50), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n757), .A2(G58), .B1(G132), .B2(new_n747), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(new_n377), .C2(new_n744), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT104), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n753), .A2(G150), .B1(G159), .B2(new_n763), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  INV_X1    g0629(.A(new_n759), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n737), .C2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  NOR2_X1   g0633(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n735), .B1(new_n823), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n735), .A2(new_n812), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n314), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n813), .A2(new_n814), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n811), .A2(new_n838), .ZN(G384));
  AND2_X1   g0639(.A1(new_n644), .A2(new_n692), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n661), .B1(new_n840), .B2(new_n691), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n695), .B1(new_n841), .B2(new_n685), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(new_n451), .B1(new_n636), .B2(new_n641), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT106), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n434), .A2(new_n445), .A3(new_n672), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n408), .B1(KEYINPUT16), .B2(new_n407), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(new_n392), .B1(new_n354), .B2(new_n659), .ZN(new_n848));
  INV_X1    g0648(.A(new_n403), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT37), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  INV_X1    g0651(.A(new_n659), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n393), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n398), .A2(new_n851), .A3(new_n403), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n399), .A2(new_n397), .A3(new_n405), .A4(new_n410), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n659), .B1(new_n847), .B2(new_n392), .ZN(new_n856));
  AOI221_X4 g0656(.A(new_n846), .B1(new_n850), .B2(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n850), .A2(new_n854), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT39), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n403), .B1(new_n409), .B2(new_n659), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n409), .A2(new_n354), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n854), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n411), .B2(new_n634), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n846), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n859), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n845), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n857), .A2(new_n860), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n808), .A2(new_n798), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n445), .A2(new_n661), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n449), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n626), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n845), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n872), .A2(new_n879), .B1(new_n634), .B2(new_n852), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n844), .B(new_n881), .ZN(new_n882));
  NOR4_X1   g0682(.A1(new_n620), .A2(new_n483), .A3(new_n526), .A4(new_n661), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n807), .B(new_n878), .C1(new_n883), .C2(new_n717), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n858), .A2(new_n859), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n846), .ZN(new_n886));
  AOI211_X1 g0686(.A(KEYINPUT40), .B(new_n884), .C1(new_n886), .C2(new_n868), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n867), .A2(new_n868), .ZN(new_n889));
  INV_X1    g0689(.A(new_n884), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(G330), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n717), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n719), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n451), .A2(G330), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n888), .B1(new_n857), .B2(new_n860), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n884), .B1(new_n868), .B2(new_n867), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n897), .A2(new_n884), .B1(new_n898), .B2(new_n888), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n451), .A3(new_n894), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n882), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n264), .B2(new_n655), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n535), .A2(new_n536), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT35), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n224), .B(new_n225), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(G116), .C1(new_n905), .C2(new_n904), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  OAI21_X1  g0708(.A(G77), .B1(new_n738), .B2(new_n377), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(new_n223), .B1(G50), .B2(new_n377), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(G1), .A3(new_n654), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n908), .A3(new_n911), .ZN(G367));
  INV_X1    g0712(.A(new_n673), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n665), .B(new_n913), .C1(new_n670), .C2(G330), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n674), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n662), .B1(new_n665), .B2(new_n913), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n539), .A2(new_n661), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n643), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n645), .A2(new_n661), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT45), .Z(new_n922));
  NAND3_X1  g0722(.A1(new_n670), .A2(G330), .A3(new_n665), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n916), .A2(new_n920), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT44), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n723), .A2(new_n724), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT107), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n677), .B(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n730), .A2(G1), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n930), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT107), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n920), .A2(new_n665), .A3(new_n913), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT42), .Z(new_n938));
  INV_X1    g0738(.A(new_n920), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n573), .B1(new_n939), .B2(new_n520), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n672), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n605), .A2(new_n672), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n615), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n614), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n938), .A2(new_n941), .B1(KEYINPUT43), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n923), .A2(new_n939), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n936), .A2(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n774), .A2(new_n778), .B1(new_n210), .B2(new_n756), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G283), .B2(new_n763), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n474), .B2(new_n737), .C1(new_n214), .C2(new_n744), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT46), .ZN(new_n958));
  INV_X1    g0758(.A(new_n761), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n457), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n785), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G311), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n830), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n746), .A2(new_n965), .ZN(new_n966));
  NOR4_X1   g0766(.A1(new_n957), .A2(new_n962), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n744), .A2(new_n314), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n761), .A2(G58), .B1(G137), .B2(new_n747), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n736), .A2(G150), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G68), .A2(new_n757), .B1(new_n753), .B2(G159), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n759), .A2(G143), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n968), .B(new_n974), .C1(G50), .C2(new_n763), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n967), .B1(new_n975), .B2(new_n271), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n735), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n943), .A2(new_n733), .A3(new_n944), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n782), .B1(new_n228), .B2(new_n312), .C1(new_n786), .C2(new_n239), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT108), .Z(new_n981));
  NAND4_X1  g0781(.A1(new_n978), .A2(new_n814), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n954), .A2(new_n982), .ZN(G387));
  NOR2_X1   g0783(.A1(new_n236), .A2(new_n468), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(new_n786), .B1(new_n680), .B2(new_n788), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n249), .A2(G50), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT50), .ZN(new_n987));
  AOI21_X1  g0787(.A(G45), .B1(G68), .B2(G77), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n680), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(G107), .B2(new_n228), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n666), .A2(new_n733), .B1(new_n782), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n785), .B1(G150), .B2(new_n747), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n753), .A2(new_n388), .B1(G50), .B2(new_n736), .ZN(new_n994));
  INV_X1    g0794(.A(G159), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n830), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n761), .A2(G77), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n608), .B2(new_n756), .C1(new_n744), .C2(new_n214), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(G68), .C2(new_n763), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n761), .A2(G294), .B1(G283), .B2(new_n757), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n737), .A2(new_n965), .B1(new_n474), .B2(new_n762), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT110), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n963), .B2(new_n774), .C1(new_n768), .C2(new_n830), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT111), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1003), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(KEYINPUT48), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n744), .A2(new_n457), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n784), .B(new_n1012), .C1(G326), .C2(new_n747), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n999), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n735), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n814), .B(new_n992), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT113), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n725), .A2(new_n915), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n725), .A2(new_n915), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n677), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n915), .A2(new_n932), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(G393));
  INV_X1    g0823(.A(new_n926), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n923), .B1(new_n922), .B2(new_n925), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n725), .A2(new_n926), .A3(new_n915), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n677), .A3(new_n1027), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n933), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n759), .A2(G150), .B1(G159), .B2(new_n736), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n819), .B1(KEYINPUT51), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n785), .B(new_n1031), .C1(G50), .C2(new_n753), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n757), .A2(G77), .B1(new_n388), .B2(new_n763), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n959), .B2(new_n377), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT51), .B2(new_n1030), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1032), .B(new_n1035), .C1(new_n831), .C2(new_n746), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n293), .B1(new_n762), .B2(new_n778), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n744), .A2(new_n210), .B1(new_n768), .B2(new_n746), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(G116), .C2(new_n757), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n816), .B2(new_n959), .C1(new_n474), .C2(new_n774), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n759), .A2(G317), .B1(G311), .B2(new_n736), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1036), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n733), .A2(new_n939), .B1(new_n1043), .B2(new_n735), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n782), .B1(new_n214), .B2(new_n228), .C1(new_n786), .C2(new_n247), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n814), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT115), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1028), .A2(new_n1029), .A3(new_n1049), .ZN(G390));
  NOR2_X1   g0850(.A1(new_n884), .A2(new_n698), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT116), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n879), .A2(new_n845), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n861), .A3(new_n870), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n799), .B1(new_n841), .B2(new_n807), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n875), .A2(new_n626), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n889), .B(new_n845), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1053), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n718), .A2(new_n719), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(G330), .A3(new_n807), .A4(new_n878), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n894), .A2(G330), .A3(new_n807), .A4(new_n878), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n1052), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1055), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n932), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1070));
  OAI211_X1 g0870(.A(G330), .B(new_n807), .C1(new_n883), .C2(new_n717), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n877), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1056), .A2(new_n1062), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n873), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n716), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT95), .B1(new_n1075), .B2(new_n711), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n711), .A2(KEYINPUT95), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(G330), .B(new_n807), .C1(new_n1078), .C2(new_n883), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n877), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1074), .B1(new_n1080), .B2(new_n1064), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n895), .B(new_n843), .C1(new_n1073), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n678), .B1(new_n1070), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n451), .B1(new_n694), .B2(new_n696), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n642), .A2(new_n1084), .A3(new_n895), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n878), .B1(new_n720), .B2(new_n807), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n873), .B1(new_n1086), .B2(new_n1051), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1056), .A2(new_n1062), .A3(new_n1072), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n631), .A2(new_n633), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n405), .A2(new_n410), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n393), .B(new_n852), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n864), .A2(new_n854), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT38), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n845), .B1(new_n857), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n693), .A2(new_n672), .A3(new_n807), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1057), .B1(new_n1096), .B2(new_n798), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n869), .B1(new_n886), .B2(new_n868), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n867), .A2(new_n869), .A3(new_n868), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1101), .B2(new_n1054), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1066), .B(new_n1089), .C1(new_n1102), .C2(new_n1053), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1068), .A2(new_n1069), .B1(new_n1083), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n812), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n830), .A2(new_n1106), .B1(new_n995), .B2(new_n756), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G137), .B2(new_n753), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n293), .B1(new_n743), .B2(G50), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1109), .C1(new_n1110), .C2(new_n746), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n959), .A2(KEYINPUT53), .A3(new_n251), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT53), .B1(new_n959), .B2(new_n251), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1112), .B(new_n1113), .C1(new_n762), .C2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1111), .B(new_n1115), .C1(G132), .C2(new_n736), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n377), .A2(new_n744), .B1(new_n959), .B2(new_n594), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n769), .A2(new_n457), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n293), .B1(new_n214), .B2(new_n762), .C1(new_n756), .C2(new_n314), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n759), .A2(G283), .B1(G294), .B2(new_n747), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n210), .B2(new_n774), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n735), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n836), .A2(new_n249), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1105), .A2(new_n814), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT118), .Z(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n1126), .ZN(G378));
  NAND2_X1  g0927(.A1(new_n624), .A2(new_n640), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT119), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1128), .B(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n270), .A2(new_n852), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n812), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n743), .A2(G58), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n997), .A2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n377), .B2(new_n756), .C1(new_n210), .C2(new_n769), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n785), .A2(new_n464), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n774), .A2(new_n214), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n608), .A2(new_n762), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n457), .B2(new_n830), .C1(new_n816), .C2(new_n746), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT58), .Z(new_n1146));
  OAI211_X1 g0946(.A(new_n1141), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1147));
  INV_X1    g0947(.A(G132), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n774), .A2(new_n1148), .B1(new_n830), .B2(new_n1110), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G150), .B2(new_n757), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n736), .A2(G128), .B1(new_n763), .B2(G137), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n959), .C2(new_n1114), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT59), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n743), .A2(G159), .B1(G124), .B2(new_n747), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n260), .A3(new_n464), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1147), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n735), .B1(new_n1146), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n836), .A2(new_n202), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1137), .A2(new_n814), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n871), .A2(new_n880), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n899), .A2(G330), .A3(new_n1135), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1135), .B1(new_n899), .B2(G330), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n892), .A2(new_n1136), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n899), .A2(G330), .A3(new_n1135), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n881), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1168), .B2(new_n932), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1085), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1164), .A2(new_n1167), .B1(new_n1103), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n677), .B1(new_n1171), .B2(KEYINPUT57), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1103), .A2(new_n1170), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1168), .A2(KEYINPUT57), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1169), .B1(new_n1172), .B2(new_n1174), .ZN(G375));
  NAND2_X1  g0975(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT122), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n757), .A2(G50), .B1(G150), .B2(new_n763), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1138), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n959), .A2(new_n995), .B1(new_n829), .B2(new_n737), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n830), .A2(new_n1148), .B1(new_n1106), .B2(new_n746), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(new_n785), .A3(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1180), .B(new_n1183), .C1(new_n774), .C2(new_n1114), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n753), .A2(G116), .B1(G107), .B2(new_n763), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT121), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G97), .B2(new_n761), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n968), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n759), .A2(G294), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n769), .A2(new_n816), .B1(new_n474), .B2(new_n746), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n271), .B(new_n1190), .C1(new_n609), .C2(new_n757), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1015), .B1(new_n1184), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n731), .B(new_n1193), .C1(new_n377), .C2(new_n836), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT123), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n877), .A2(new_n812), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT120), .Z(new_n1197));
  AOI22_X1  g0997(.A1(new_n1176), .A2(new_n932), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n930), .B1(new_n1176), .B2(new_n1170), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1089), .ZN(G381));
  OR2_X1    g1000(.A1(G381), .A2(G384), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1168), .A2(new_n932), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1159), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1162), .A2(new_n1163), .A3(new_n1161), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n881), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1055), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1206), .A2(new_n1059), .A3(new_n1082), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1204), .A2(new_n1205), .B1(new_n1207), .B2(new_n1085), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n678), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1171), .A2(KEYINPUT57), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1203), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1213), .A2(new_n1126), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(G393), .A2(G396), .ZN(new_n1217));
  INV_X1    g1017(.A(G390), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n954), .A3(new_n982), .ZN(new_n1219));
  OR4_X1    g1019(.A1(new_n1201), .A2(new_n1216), .A3(new_n1217), .A4(new_n1219), .ZN(G407));
  INV_X1    g1020(.A(G213), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(G343), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT124), .B1(new_n1216), .B2(new_n1223), .ZN(new_n1224));
  OR3_X1    g1024(.A1(new_n1216), .A2(KEYINPUT124), .A3(new_n1223), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1224), .A4(new_n1225), .ZN(G409));
  NAND2_X1  g1026(.A1(new_n1171), .A2(new_n930), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1104), .A2(new_n1126), .A3(new_n1169), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1223), .B(new_n1228), .C1(new_n1212), .C2(new_n1215), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1176), .B2(new_n1170), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1085), .A2(new_n1087), .A3(KEYINPUT60), .A4(new_n1088), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n677), .A4(new_n1082), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(G384), .A3(new_n1198), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G384), .B1(new_n1233), .B2(new_n1198), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT62), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1236), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT126), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(new_n1234), .ZN(new_n1242));
  INV_X1    g1042(.A(G2897), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1223), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT126), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1244), .B1(new_n1246), .B2(new_n1242), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1229), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1222), .B1(G375), .B2(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1237), .A4(new_n1228), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1239), .A2(new_n1249), .A3(new_n1250), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT127), .B1(G387), .B2(new_n1218), .ZN(new_n1255));
  INV_X1    g1055(.A(G396), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(G393), .B(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(G390), .B1(new_n954), .B2(new_n982), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n954), .A2(G390), .A3(new_n982), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1255), .A2(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(G393), .B(G396), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1218), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n954), .A2(G390), .A3(new_n982), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(KEYINPUT127), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1254), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1237), .A4(new_n1228), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n1265), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1247), .B1(new_n1251), .B2(new_n1228), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1245), .ZN(new_n1271));
  XOR2_X1   g1071(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1274), .ZN(G405));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1216), .A2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1277), .A2(new_n1237), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1238), .B1(new_n1216), .B2(new_n1276), .ZN(new_n1279));
  OR3_X1    g1079(.A1(new_n1278), .A2(new_n1265), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1265), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(G402));
endmodule


