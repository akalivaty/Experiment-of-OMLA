//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  OAI211_X1 g002(.A(new_n187), .B(G146), .C1(new_n188), .C2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n191), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n203), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n204), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT64), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n194), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n194), .A2(KEYINPUT64), .A3(new_n216), .A4(new_n218), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n209), .B1(new_n212), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G116), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G113), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT67), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n230), .B1(new_n235), .B2(new_n229), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT28), .B1(new_n223), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT26), .B(G101), .Z(new_n239));
  NOR2_X1   g053(.A1(G237), .A2(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G210), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n239), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n209), .A2(KEYINPUT68), .B1(new_n222), .B2(new_n212), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n208), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n248), .A3(new_n236), .A4(new_n250), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n192), .A2(new_n193), .A3(new_n214), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n221), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n212), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n196), .A2(KEYINPUT68), .A3(new_n204), .A4(new_n207), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n258), .A2(new_n236), .A3(new_n250), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n235), .A2(new_n229), .ZN(new_n262));
  INV_X1    g076(.A(new_n230), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n250), .A3(new_n259), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n251), .A2(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n238), .B(new_n246), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT74), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n251), .A2(new_n261), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(new_n256), .B2(new_n257), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n220), .A2(new_n274), .A3(new_n221), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n212), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT66), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n196), .A2(new_n278), .A3(new_n204), .A4(new_n207), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n236), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n272), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n276), .A2(new_n280), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n251), .A2(new_n261), .B1(new_n284), .B2(new_n264), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n285), .B2(new_n267), .ZN(new_n286));
  INV_X1    g100(.A(new_n244), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n282), .A2(new_n286), .A3(new_n287), .A4(new_n238), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n291), .A3(new_n280), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(KEYINPUT30), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n294), .A2(new_n264), .B1(new_n251), .B2(new_n261), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(new_n287), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(new_n245), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n288), .A2(new_n289), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n271), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G472), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(G472), .A2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n286), .A3(new_n238), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n244), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT31), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n264), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n251), .A2(new_n261), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n308), .A2(new_n309), .A3(new_n287), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n295), .B2(new_n287), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n305), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n313), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n301), .ZN(new_n319));
  INV_X1    g133(.A(new_n303), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n287), .A3(new_n310), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT31), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n295), .A2(new_n308), .A3(new_n287), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n244), .B2(new_n306), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT72), .B(new_n320), .C1(new_n325), .C2(new_n305), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n300), .A2(new_n316), .A3(new_n319), .A4(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT100), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT9), .B(G234), .Z(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(G217), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT94), .B1(new_n187), .B2(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT94), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n188), .A3(G143), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT95), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n187), .A2(G128), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n198), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n335), .B1(new_n188), .B2(G143), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n187), .A2(KEYINPUT94), .A3(G128), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT95), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(G134), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G122), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT93), .B1(new_n350), .B2(G116), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n226), .A3(G122), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(G116), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n351), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n356), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n351), .B2(new_n353), .ZN(new_n361));
  OAI21_X1  g175(.A(G107), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT96), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(G107), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n349), .A2(new_n357), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT13), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n337), .B1(new_n367), .B2(new_n339), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT13), .B1(new_n187), .B2(G128), .ZN(new_n369));
  OAI21_X1  g183(.A(G134), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n354), .A2(new_n356), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G107), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n357), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n342), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n329), .B(new_n333), .C1(new_n366), .C2(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n340), .A2(new_n341), .A3(new_n198), .ZN(new_n376));
  AOI21_X1  g190(.A(G134), .B1(new_n346), .B2(new_n347), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n357), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n363), .A2(new_n365), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT98), .B1(new_n380), .B2(new_n332), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n380), .B2(new_n332), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n366), .A2(KEYINPUT97), .A3(new_n374), .A4(new_n333), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n269), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n384), .B(new_n385), .C1(new_n375), .C2(new_n381), .ZN(new_n391));
  INV_X1    g205(.A(new_n389), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n269), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(G234), .A2(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(G952), .A3(new_n331), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT99), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT21), .B(G898), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(G902), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n397), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n406), .B(KEYINPUT90), .Z(new_n407));
  NAND3_X1  g221(.A1(new_n240), .A2(G143), .A3(G214), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(G143), .B1(new_n240), .B2(G214), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n240), .A2(G214), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n187), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n202), .A3(new_n408), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n417));
  INV_X1    g231(.A(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G125), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n417), .B(G146), .C1(KEYINPUT16), .C2(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(G125), .B(G140), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT19), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n424), .A3(new_n190), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n416), .B(new_n190), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n413), .B(new_n408), .C1(new_n428), .C2(new_n202), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n427), .B(new_n429), .C1(new_n428), .C2(new_n411), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT89), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  INV_X1    g247(.A(G104), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n426), .A2(new_n430), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n411), .A2(new_n414), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n417), .B1(KEYINPUT16), .B2(new_n419), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n190), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT17), .B(G131), .C1(new_n409), .C2(new_n410), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n420), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n435), .A3(new_n430), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n407), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n405), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n445), .A2(new_n435), .A3(new_n430), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n435), .B1(new_n431), .B2(KEYINPUT89), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n438), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n452), .C2(new_n407), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n448), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n435), .B1(new_n445), .B2(new_n430), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n269), .B1(new_n450), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT92), .B(G475), .Z(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n328), .B1(new_n404), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n391), .A2(new_n269), .A3(new_n392), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n392), .B1(new_n391), .B2(new_n269), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n455), .A2(new_n459), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT100), .A4(new_n403), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G221), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n330), .B2(new_n269), .ZN(new_n469));
  INV_X1    g283(.A(G469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n355), .A2(G104), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n434), .A2(G107), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n475));
  OAI211_X1 g289(.A(G104), .B(new_n355), .C1(new_n475), .C2(KEYINPUT80), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n477));
  INV_X1    g291(.A(new_n471), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n476), .B(new_n472), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n196), .B(new_n474), .C1(new_n479), .C2(G101), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT10), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT3), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n471), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G101), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n476), .A4(new_n472), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n196), .A4(new_n474), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n212), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n479), .A2(G101), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT4), .A3(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n479), .A2(new_n494), .A3(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n222), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT81), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT81), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n490), .A2(new_n496), .A3(new_n499), .A4(new_n491), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(G110), .B(G140), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n331), .A2(G227), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n487), .A2(new_n474), .ZN(new_n505));
  INV_X1    g319(.A(new_n196), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n480), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n501), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n490), .A2(new_n496), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n212), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n504), .B1(new_n501), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n470), .B(new_n269), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n501), .A2(new_n504), .A3(new_n513), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n498), .A2(new_n500), .B1(new_n212), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n504), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n470), .A4(new_n269), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n501), .A2(new_n516), .A3(new_n504), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n501), .A2(new_n513), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n504), .B1(new_n527), .B2(KEYINPUT83), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT83), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n501), .A2(new_n529), .A3(new_n513), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G469), .B1(new_n531), .B2(G902), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n469), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(G110), .B(G122), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n505), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT5), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n224), .A3(G116), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(G113), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n235), .B2(new_n537), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n263), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n264), .A2(new_n493), .A3(new_n495), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(KEYINPUT6), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n542), .A3(new_n535), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT86), .A4(new_n535), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n220), .A2(G125), .A3(new_n221), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n196), .A2(G125), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n331), .A2(G224), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT88), .Z(new_n560));
  OAI21_X1  g374(.A(new_n539), .B1(new_n537), .B2(new_n228), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n536), .A2(new_n263), .A3(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n540), .A2(new_n263), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n505), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n534), .B(KEYINPUT8), .Z(new_n568));
  NAND2_X1  g382(.A1(new_n555), .A2(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n552), .A2(new_n553), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n554), .A2(KEYINPUT7), .A3(new_n555), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n567), .A2(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n547), .A2(new_n548), .ZN(new_n573));
  AOI21_X1  g387(.A(G902), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n558), .A2(new_n560), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n560), .B1(new_n558), .B2(new_n574), .ZN(new_n576));
  OAI21_X1  g390(.A(G214), .B1(G237), .B2(G902), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT85), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n467), .A2(new_n533), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n443), .A2(new_n420), .ZN(new_n581));
  XOR2_X1   g395(.A(KEYINPUT24), .B(G110), .Z(new_n582));
  XNOR2_X1  g396(.A(G119), .B(G128), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT23), .B1(new_n188), .B2(G119), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n188), .A2(G119), .ZN(new_n586));
  MUX2_X1   g400(.A(KEYINPUT23), .B(new_n585), .S(new_n586), .Z(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G110), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n581), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OAI22_X1  g403(.A1(new_n587), .A2(G110), .B1(new_n583), .B2(new_n582), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n590), .B(new_n420), .C1(G146), .C2(new_n421), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT22), .B(G137), .ZN(new_n593));
  INV_X1    g407(.A(G234), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n468), .A2(new_n594), .A3(G953), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n593), .B(new_n595), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n589), .A2(new_n591), .A3(new_n596), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n269), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT25), .ZN(new_n601));
  OAI21_X1  g415(.A(G217), .B1(new_n594), .B2(G902), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT76), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT77), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT25), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n598), .A2(new_n605), .A3(new_n269), .A4(new_n599), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n598), .A2(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n269), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n609), .B(KEYINPUT78), .Z(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n327), .A2(new_n580), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND2_X1  g432(.A1(new_n525), .A2(new_n532), .ZN(new_n619));
  INV_X1    g433(.A(new_n469), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n317), .A2(new_n304), .ZN(new_n622));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n307), .B2(new_n313), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n622), .B(new_n616), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT101), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n579), .A2(new_n403), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n382), .B2(new_n386), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n380), .A2(new_n332), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n366), .A2(new_n374), .A3(new_n333), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(KEYINPUT33), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n630), .A2(G478), .A3(new_n269), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n387), .A2(new_n388), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n460), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n627), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n628), .ZN(new_n642));
  INV_X1    g456(.A(new_n464), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n454), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n447), .A2(KEYINPUT102), .A3(new_n448), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n449), .A3(new_n453), .A4(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n459), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n642), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NAND2_X1  g467(.A1(new_n317), .A2(new_n269), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n314), .B1(new_n654), .B2(G472), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n597), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n592), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n610), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n607), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n580), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  OAI21_X1  g476(.A(new_n396), .B1(G900), .B2(new_n400), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n647), .A2(new_n459), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n464), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n533), .A2(new_n579), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n327), .A2(new_n659), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT103), .B(G128), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G30));
  XOR2_X1   g483(.A(new_n663), .B(KEYINPUT39), .Z(new_n670));
  NOR2_X1   g484(.A1(new_n621), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  NOR2_X1   g486(.A1(new_n575), .A2(new_n576), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT38), .Z(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n464), .A2(new_n465), .ZN(new_n676));
  INV_X1    g490(.A(new_n578), .ZN(new_n677));
  INV_X1    g491(.A(new_n659), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT104), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n266), .A2(new_n287), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n287), .B2(new_n295), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n682), .B2(G902), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n319), .A2(new_n326), .A3(new_n316), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n675), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n672), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n187), .ZN(G45));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n677), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n621), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n636), .A2(new_n460), .A3(new_n663), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n327), .A2(new_n689), .A3(new_n659), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  AOI21_X1  g507(.A(new_n470), .B1(new_n523), .B2(new_n269), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n469), .B(new_n694), .C1(new_n520), .C2(new_n524), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n319), .A2(new_n326), .A3(new_n316), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT29), .B1(new_n288), .B2(new_n289), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n296), .C1(new_n289), .C2(new_n288), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n623), .B1(new_n698), .B2(new_n271), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n616), .B(new_n695), .C1(new_n696), .C2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n638), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  INV_X1    g520(.A(new_n700), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n650), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n700), .A2(KEYINPUT106), .A3(new_n649), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT107), .B(G116), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  AOI21_X1  g526(.A(new_n694), .B1(new_n520), .B2(new_n524), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n620), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n688), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n467), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n327), .A4(new_n659), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n659), .B1(new_n696), .B2(new_n699), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n467), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT108), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT109), .B(G119), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G21));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n265), .A2(new_n264), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n310), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT28), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n287), .B1(new_n728), .B2(new_n238), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n729), .B2(new_n312), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n267), .B1(new_n310), .B2(new_n726), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n244), .B1(new_n731), .B2(new_n237), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n322), .A2(new_n732), .A3(KEYINPUT110), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n323), .A3(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n654), .A2(G472), .B1(new_n734), .B2(new_n304), .ZN(new_n735));
  INV_X1    g549(.A(new_n612), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n695), .A2(new_n676), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n628), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n350), .ZN(G24));
  AND4_X1   g554(.A1(KEYINPUT111), .A2(new_n636), .A3(new_n460), .A4(new_n663), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n634), .A2(new_n635), .B1(new_n455), .B2(new_n459), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n743), .B2(new_n663), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n735), .A2(new_n659), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n747), .A3(new_n715), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND2_X1  g563(.A1(new_n622), .A2(new_n302), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n751), .A2(new_n317), .A3(KEYINPUT32), .A4(new_n304), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n314), .B2(KEYINPUT32), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n736), .B1(new_n754), .B2(new_n699), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n558), .A2(new_n574), .ZN(new_n756));
  INV_X1    g570(.A(new_n560), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n558), .A2(new_n560), .A3(new_n574), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n578), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n619), .A2(new_n760), .A3(new_n620), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n744), .B2(new_n741), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT42), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n533), .A2(new_n760), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n742), .B2(new_n745), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n327), .A4(new_n616), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n202), .ZN(G33));
  INV_X1    g583(.A(new_n616), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n319), .A2(new_n316), .A3(new_n326), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n300), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n665), .A4(new_n761), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n761), .B(new_n616), .C1(new_n696), .C2(new_n699), .ZN(new_n775));
  INV_X1    g589(.A(new_n665), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT113), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  XOR2_X1   g593(.A(new_n531), .B(KEYINPUT45), .Z(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(G469), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n525), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n620), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(new_n670), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n760), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n460), .B1(new_n634), .B2(new_n635), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT43), .Z(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(new_n655), .A3(new_n678), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  NAND2_X1  g611(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n327), .A2(new_n616), .A3(new_n789), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n800), .B(new_n620), .C1(new_n784), .C2(new_n785), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n798), .A2(new_n691), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  INV_X1    g617(.A(new_n713), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT115), .Z(new_n806));
  NAND4_X1  g620(.A1(new_n790), .A2(new_n736), .A3(new_n620), .A4(new_n677), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT114), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n684), .B1(KEYINPUT49), .B2(new_n804), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(new_n808), .A3(new_n674), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n791), .A2(new_n396), .A3(new_n737), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n760), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n798), .A2(new_n801), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n713), .A2(new_n469), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n578), .A3(new_n674), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT50), .B1(new_n816), .B2(new_n714), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n695), .A2(new_n760), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n684), .A2(new_n818), .A3(new_n770), .A4(new_n396), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n465), .A3(new_n635), .A4(new_n634), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n791), .A2(new_n396), .A3(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n747), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n816), .A2(KEYINPUT50), .A3(new_n714), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n815), .A2(new_n823), .A3(new_n828), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n318), .A2(KEYINPUT112), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n314), .A2(new_n751), .A3(KEYINPUT32), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n830), .A2(new_n831), .B1(new_n302), .B2(new_n622), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n612), .B1(new_n832), .B2(new_n300), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n821), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT121), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT48), .ZN(new_n836));
  OAI211_X1 g650(.A(G952), .B(new_n331), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n827), .A2(new_n829), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n819), .A2(new_n743), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n834), .A2(KEYINPUT121), .A3(KEYINPUT48), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n811), .A2(new_n715), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT120), .Z(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n462), .A2(new_n463), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT116), .B1(new_n390), .B2(new_n393), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n465), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT117), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n465), .C1(new_n847), .C2(new_n848), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n637), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n642), .A3(new_n626), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n617), .A2(new_n660), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n761), .A2(new_n659), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n746), .A2(new_n735), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n847), .A2(new_n848), .A3(new_n664), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n696), .B2(new_n699), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n768), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n737), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n642), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n863), .A2(new_n738), .B1(new_n700), .B2(new_n701), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n718), .B2(new_n721), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(new_n710), .A3(new_n778), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n679), .ZN(new_n867));
  INV_X1    g681(.A(new_n663), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n469), .B(new_n868), .C1(new_n525), .C2(new_n532), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n684), .A2(new_n673), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n621), .A2(new_n679), .A3(new_n868), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n673), .A4(new_n684), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n692), .A2(new_n667), .A3(new_n748), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT52), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n692), .A2(new_n667), .A3(new_n748), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n874), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n845), .B1(new_n866), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n855), .A2(new_n860), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n833), .A2(new_n765), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n766), .B(new_n616), .C1(new_n696), .C2(new_n699), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n885), .A2(KEYINPUT42), .B1(new_n887), .B2(new_n765), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n888), .A3(new_n778), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n702), .A2(new_n739), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n722), .C1(new_n708), .C2(new_n709), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n735), .A2(new_n579), .A3(new_n659), .A4(new_n695), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n741), .A2(new_n744), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n678), .B1(new_n771), .B2(new_n300), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n896), .B2(new_n666), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n879), .A2(new_n880), .A3(new_n897), .A4(new_n692), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n892), .A2(new_n900), .A3(KEYINPUT53), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n883), .A2(KEYINPUT54), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT54), .B1(new_n883), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n844), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n902), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n843), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(G952), .A2(G953), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n810), .B1(new_n908), .B2(new_n909), .ZN(G75));
  AOI21_X1  g724(.A(new_n269), .B1(new_n883), .B2(new_n901), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n560), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n551), .B(new_n556), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n331), .A2(G952), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G51));
  NAND3_X1  g733(.A1(new_n911), .A2(G469), .A3(new_n780), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n782), .A2(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n906), .A2(new_n902), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n782), .A2(KEYINPUT57), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n523), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n918), .B1(new_n921), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n452), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n452), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n918), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n630), .A2(new_n633), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT123), .Z(new_n934));
  NOR4_X1   g748(.A1(new_n903), .A2(new_n904), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n932), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n905), .A2(new_n907), .A3(new_n936), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n918), .B(new_n935), .C1(new_n937), .C2(new_n934), .ZN(G63));
  NAND2_X1  g752(.A1(new_n883), .A2(new_n901), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT124), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n944), .B(new_n941), .C1(new_n883), .C2(new_n901), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n657), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n866), .A2(new_n845), .A3(new_n882), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT53), .B1(new_n892), .B2(new_n900), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n944), .ZN(new_n950));
  INV_X1    g764(.A(new_n608), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n939), .A2(KEYINPUT124), .A3(new_n942), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n918), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n946), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n946), .A2(new_n953), .A3(KEYINPUT61), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(G66));
  AOI21_X1  g773(.A(new_n331), .B1(new_n398), .B2(G224), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n891), .A2(new_n855), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n964), .B2(new_n331), .ZN(new_n965));
  INV_X1    g779(.A(new_n551), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G898), .B2(new_n331), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n965), .B(new_n967), .Z(G69));
  AOI21_X1  g782(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND2_X1  g786(.A1(G900), .A2(G953), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n294), .B(KEYINPUT126), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n422), .A2(new_n424), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(new_n976));
  AND3_X1   g790(.A1(new_n796), .A2(new_n888), .A3(new_n802), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n787), .A2(new_n575), .A3(new_n576), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(new_n677), .A3(new_n676), .A4(new_n833), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n977), .A2(new_n778), .A3(new_n878), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n973), .B(new_n976), .C1(new_n980), .C2(G953), .ZN(new_n981));
  INV_X1    g795(.A(new_n976), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n775), .A2(new_n670), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n853), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n796), .A2(new_n802), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n878), .B1(new_n685), .B2(new_n672), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT62), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n982), .B1(new_n988), .B2(G953), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n971), .B(new_n972), .C1(new_n981), .C2(new_n989), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n970), .A2(new_n981), .A3(new_n969), .A4(new_n989), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G72));
  NAND3_X1  g806(.A1(new_n988), .A2(new_n963), .A3(new_n962), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  AOI21_X1  g809(.A(new_n295), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n918), .B1(new_n996), .B2(new_n287), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n995), .B1(new_n980), .B2(new_n964), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n244), .A3(new_n295), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n296), .A2(new_n321), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n939), .A2(new_n995), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(G57));
endmodule


