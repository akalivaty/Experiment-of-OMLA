//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(new_n204), .ZN(new_n214));
  AND2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT74), .B1(new_n215), .B2(new_n211), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n210), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n205), .B1(new_n215), .B2(new_n211), .ZN(new_n218));
  INV_X1    g017(.A(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(G148gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n218), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT76), .B1(new_n217), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n219), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n204), .B1(new_n212), .B2(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n214), .A3(new_n216), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT76), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n225), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n228), .A2(new_n229), .A3(new_n236), .A4(new_n238), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n203), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n225), .A2(KEYINPUT3), .A3(new_n231), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n236), .A2(new_n238), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n217), .A2(new_n224), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n241), .B(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n243), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n203), .A4(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT0), .ZN(new_n258));
  XNOR2_X1  g057(.A(G57gat), .B(G85gat), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT6), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n260), .A3(new_n255), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n254), .B2(new_n255), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT6), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT23), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT24), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(G183gat), .A3(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n270), .A2(new_n272), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n280), .A2(KEYINPUT24), .A3(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n268), .B(KEYINPUT25), .C1(new_n277), .C2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n270), .A2(new_n276), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n272), .A2(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n268), .A2(KEYINPUT25), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(KEYINPUT24), .A3(new_n281), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(KEYINPUT66), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(new_n269), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n302), .A3(new_n291), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n296), .A2(new_n299), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n307), .A3(new_n279), .ZN(new_n308));
  NAND2_X1  g107(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n308), .A2(new_n310), .B1(G183gat), .B2(G190gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n312), .A2(new_n279), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n304), .A2(new_n311), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n289), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n289), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n315), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n319), .A2(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT71), .B(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G197gat), .B(G204gat), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n329), .B2(new_n331), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(KEYINPUT72), .B(new_n320), .C1(new_n319), .C2(KEYINPUT29), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n308), .A2(new_n310), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n314), .A2(new_n339), .A3(new_n281), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n317), .B1(new_n340), .B2(new_n304), .ZN(new_n341));
  INV_X1    g140(.A(new_n318), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n322), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n321), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n315), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n321), .B1(new_n346), .B2(new_n289), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n338), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n337), .B1(new_n350), .B2(new_n336), .ZN(new_n351));
  XOR2_X1   g150(.A(G8gat), .B(G36gat), .Z(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT73), .ZN(new_n353));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n265), .A2(new_n267), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT38), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n320), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n348), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n336), .B1(new_n360), .B2(new_n338), .ZN(new_n361));
  INV_X1    g160(.A(new_n336), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT37), .B1(new_n325), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n355), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n360), .B2(new_n338), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n337), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(KEYINPUT37), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n202), .B1(new_n357), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT37), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n355), .B1(new_n351), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n263), .B(new_n260), .C1(new_n254), .C2(new_n255), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n266), .A2(KEYINPUT6), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n264), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT86), .A4(new_n356), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n372), .B1(new_n371), .B2(new_n351), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT38), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n228), .A2(new_n229), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n344), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n336), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n344), .B1(new_n334), .B2(new_n335), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n332), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT71), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G211gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT22), .B1(new_n395), .B2(G218gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n396), .B2(new_n330), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n397), .B2(new_n333), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n249), .B1(new_n398), .B2(KEYINPUT80), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n383), .B1(new_n389), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n386), .B1(new_n400), .B2(KEYINPUT81), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT3), .B1(new_n387), .B2(new_n388), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(KEYINPUT80), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n248), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n401), .A2(new_n406), .B1(G228gat), .B2(G233gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n384), .B2(new_n336), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n225), .B(new_n231), .C1(new_n398), .C2(KEYINPUT3), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(G22gat), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n385), .B1(new_n404), .B2(new_n405), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT81), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n422), .A3(KEYINPUT83), .ZN(new_n423));
  XOR2_X1   g222(.A(G78gat), .B(G106gat), .Z(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(G22gat), .C1(new_n407), .C2(new_n413), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n406), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n431), .A2(new_n408), .B1(new_n419), .B2(new_n420), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n426), .B1(new_n432), .B2(new_n418), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(G22gat), .C1(new_n407), .C2(new_n413), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT39), .B1(new_n242), .B2(new_n244), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n261), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n262), .B1(new_n442), .B2(KEYINPUT40), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(KEYINPUT40), .A3(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n444), .A2(new_n445), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n356), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n351), .A2(KEYINPUT30), .A3(new_n355), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n367), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n429), .A2(new_n436), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n382), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G227gat), .ZN(new_n455));
  INV_X1    g254(.A(G233gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n343), .A2(new_n239), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n319), .A2(new_n247), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT32), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G43gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n319), .A2(new_n247), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n239), .B(new_n289), .C1(new_n316), .C2(new_n318), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT70), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n472), .A3(KEYINPUT32), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n463), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n469), .B(KEYINPUT32), .C1(new_n470), .C2(new_n466), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n467), .A2(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n458), .ZN(new_n479));
  NOR4_X1   g278(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT34), .A4(new_n457), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(new_n481), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT36), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n265), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n264), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n267), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n451), .A2(new_n367), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT30), .B1(new_n351), .B2(new_n355), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n429), .A2(new_n436), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n486), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n485), .B1(new_n429), .B2(new_n436), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n429), .A2(new_n436), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n483), .A2(new_n484), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n452), .A2(KEYINPUT35), .A3(new_n377), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n454), .A2(new_n500), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  OR2_X1    g309(.A1(G43gat), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G43gat), .A2(G50gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n517), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n513), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n513), .B1(G29gat), .B2(G36gat), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT88), .B(G50gat), .Z(new_n526));
  OAI211_X1 g325(.A(new_n510), .B(new_n512), .C1(new_n526), .C2(G43gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n527), .A3(new_n518), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT90), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(KEYINPUT17), .A3(new_n528), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT91), .Z(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G1gat), .B2(new_n535), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n532), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n529), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n540), .B(new_n529), .Z(new_n547));
  XOR2_X1   g346(.A(new_n542), .B(KEYINPUT13), .Z(new_n548));
  AOI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n541), .A2(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n542), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT11), .B(G169gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT12), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n549), .B2(new_n551), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n509), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT93), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(KEYINPUT95), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(KEYINPUT95), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G85gat), .B2(G92gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n582), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(KEYINPUT97), .A3(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n534), .A3(new_n532), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT98), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n529), .A3(new_n587), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n591), .A2(KEYINPUT98), .B1(KEYINPUT41), .B2(new_n564), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n592), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n589), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n569), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n592), .B1(new_n590), .B2(new_n595), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n597), .A3(new_n589), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n568), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G71gat), .B(G78gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n586), .A2(new_n587), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n584), .A2(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n581), .A2(new_n611), .A3(new_n583), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n605), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n605), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT100), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n620), .A2(new_n628), .A3(new_n622), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n620), .A2(new_n622), .ZN(new_n630));
  INV_X1    g429(.A(new_n625), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n627), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G127gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n540), .B1(new_n633), .B2(new_n611), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n640), .B(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n604), .A2(new_n632), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n562), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n490), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n493), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT101), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(G8gat), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT16), .B(G8gat), .Z(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(KEYINPUT42), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n652), .B(new_n654), .C1(new_n656), .C2(KEYINPUT42), .ZN(G1325gat));
  XNOR2_X1  g456(.A(new_n505), .B(KEYINPUT36), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n647), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n485), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n647), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n647), .A2(new_n504), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n629), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n630), .A2(new_n631), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n645), .ZN(new_n668));
  INV_X1    g467(.A(new_n604), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT102), .Z(new_n671));
  NAND2_X1  g470(.A1(new_n562), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(G29gat), .A3(new_n490), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT45), .Z(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n509), .B2(new_n604), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n493), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT79), .B1(new_n490), .B2(new_n493), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n499), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n454), .A2(new_n679), .A3(new_n658), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT35), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n501), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n683), .B2(new_n507), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n669), .ZN(new_n685));
  INV_X1    g484(.A(new_n560), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(KEYINPUT103), .A3(new_n558), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n559), .B2(new_n560), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n685), .A3(new_n691), .A4(new_n668), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n490), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n693), .ZN(G1328gat));
  NOR3_X1   g493(.A1(new_n672), .A2(G36gat), .A3(new_n493), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n692), .B2(new_n493), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  NOR2_X1   g497(.A1(new_n672), .A2(new_n485), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n486), .A2(G43gat), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n699), .A2(G43gat), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g501(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n499), .A2(new_n526), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n672), .A2(new_n504), .ZN(new_n705));
  OAI221_X1 g504(.A(new_n703), .B1(new_n692), .B2(new_n704), .C1(new_n705), .C2(new_n526), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT104), .A2(KEYINPUT48), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n706), .B(new_n707), .Z(G1331gat));
  INV_X1    g507(.A(new_n645), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n691), .A2(new_n709), .A3(new_n669), .A4(new_n632), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n684), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n490), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g513(.A(new_n493), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT105), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  INV_X1    g518(.A(new_n711), .ZN(new_n720));
  OAI21_X1  g519(.A(G71gat), .B1(new_n720), .B2(new_n658), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n485), .A2(G71gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g523(.A1(new_n711), .A2(new_n499), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT106), .B(G78gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n509), .A2(new_n604), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n691), .A2(new_n645), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n729), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n669), .A4(new_n730), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n454), .A2(new_n679), .A3(new_n658), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n507), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n669), .B(new_n730), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n632), .ZN(new_n742));
  INV_X1    g541(.A(G85gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n743), .A3(new_n712), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n691), .A2(new_n645), .A3(new_n632), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n676), .A2(new_n685), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n490), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  OAI21_X1  g549(.A(G92gat), .B1(new_n747), .B2(new_n493), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n632), .A2(G92gat), .A3(new_n493), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n740), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n740), .B2(new_n753), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n750), .B(new_n751), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n732), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n753), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n759), .B2(new_n750), .ZN(G1337gat));
  AOI21_X1  g559(.A(G99gat), .B1(new_n742), .B2(new_n505), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n486), .A2(G99gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n746), .B2(new_n762), .ZN(G1338gat));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n676), .A2(new_n499), .A3(new_n685), .A4(new_n745), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(G106gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n632), .A2(new_n504), .A3(G106gat), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT111), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770));
  INV_X1    g569(.A(new_n768), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n770), .B(new_n771), .C1(new_n739), .C2(new_n732), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n767), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n766), .A2(new_n765), .A3(G106gat), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n764), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n766), .B2(KEYINPUT112), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(KEYINPUT112), .B2(new_n766), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n740), .B2(new_n768), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT113), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n769), .A2(new_n772), .ZN(new_n782));
  INV_X1    g581(.A(new_n767), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n783), .A3(new_n774), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n779), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n604), .A2(new_n632), .A3(new_n645), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n691), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n646), .A2(KEYINPUT114), .A3(new_n690), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n550), .A2(new_n542), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n547), .A2(new_n548), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n555), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n558), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n667), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n618), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n611), .B1(new_n581), .B2(new_n583), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n615), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n586), .A2(new_n587), .A3(new_n613), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n621), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n620), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n621), .B1(new_n802), .B2(new_n803), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n625), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT55), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n665), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n799), .B1(new_n690), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n604), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n669), .A2(new_n798), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n794), .B1(new_n818), .B2(new_n709), .ZN(new_n819));
  INV_X1    g618(.A(new_n501), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n490), .A2(new_n452), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n561), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n690), .A2(G113gat), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n824), .B2(new_n827), .ZN(G1340gat));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n667), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n645), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n637), .A2(KEYINPUT116), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n604), .A2(new_n490), .A3(new_n452), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n821), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n824), .B2(new_n604), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n792), .A2(new_n793), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n805), .A2(new_n808), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n842), .A2(KEYINPUT55), .B1(new_n627), .B2(new_n629), .ZN(new_n843));
  INV_X1    g642(.A(new_n561), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n811), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n669), .B1(new_n845), .B2(new_n799), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n816), .A2(new_n813), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n709), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n840), .B(new_n504), .C1(new_n841), .C2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n819), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n499), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n840), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n658), .A2(new_n822), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n854), .A2(new_n691), .B1(new_n220), .B2(new_n222), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n851), .A2(new_n853), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n561), .A2(G141gat), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT117), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(KEYINPUT58), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n220), .A2(new_n222), .ZN(new_n862));
  INV_X1    g661(.A(new_n853), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n819), .A2(new_n504), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n849), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n866), .B2(new_n561), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n860), .A2(new_n868), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n856), .A2(new_n208), .A3(new_n667), .ZN(new_n870));
  AOI211_X1 g669(.A(KEYINPUT59), .B(new_n208), .C1(new_n854), .C2(new_n667), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n504), .A2(new_n840), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n646), .A2(new_n561), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n848), .B2(new_n876), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n878), .A2(new_n879), .A3(new_n504), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n667), .A3(new_n863), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n872), .B1(new_n882), .B2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n870), .B1(new_n871), .B2(new_n883), .ZN(G1345gat));
  OAI21_X1  g683(.A(G155gat), .B1(new_n866), .B2(new_n709), .ZN(new_n885));
  INV_X1    g684(.A(G155gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n856), .A2(new_n886), .A3(new_n645), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(new_n887), .A3(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n866), .B2(new_n604), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n486), .A2(G162gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n864), .A2(new_n835), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n712), .A2(new_n493), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n505), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n504), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n900), .B2(new_n899), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n850), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n293), .A3(new_n561), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n843), .A2(new_n689), .A3(new_n687), .A4(new_n811), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n669), .B1(new_n905), .B2(new_n799), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n709), .B1(new_n906), .B2(new_n847), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n712), .B1(new_n907), .B2(new_n841), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n452), .B1(new_n908), .B2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n910), .B(new_n712), .C1(new_n907), .C2(new_n841), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n909), .A2(new_n820), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n691), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n904), .B1(new_n913), .B2(new_n293), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n903), .B2(new_n632), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n910), .B1(new_n819), .B2(new_n712), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n452), .A4(new_n501), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n667), .A2(new_n294), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1349gat));
  OAI21_X1  g719(.A(G183gat), .B1(new_n903), .B2(new_n709), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n645), .A2(new_n312), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT123), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n918), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n921), .C1(new_n924), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n903), .B2(new_n604), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n669), .A2(new_n279), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n918), .B2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n909), .A2(new_n911), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n486), .A2(new_n504), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT124), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n691), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(G197gat), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n658), .A2(new_n898), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT125), .Z(new_n945));
  AND2_X1   g744(.A1(new_n881), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n561), .A2(new_n943), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n942), .A2(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND2_X1  g747(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n632), .A2(G204gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n936), .A2(new_n937), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n952));
  INV_X1    g751(.A(new_n950), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n938), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n879), .A2(new_n504), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT57), .B1(new_n955), .B2(new_n877), .ZN(new_n956));
  INV_X1    g755(.A(new_n874), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n667), .B(new_n945), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n958), .A2(KEYINPUT127), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n951), .B(new_n954), .C1(new_n960), .C2(new_n961), .ZN(G1353gat));
  NAND4_X1  g761(.A1(new_n939), .A2(new_n327), .A3(new_n645), .A4(new_n941), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n881), .A2(new_n645), .A3(new_n945), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  NAND4_X1  g766(.A1(new_n939), .A2(new_n328), .A3(new_n669), .A4(new_n941), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n946), .A2(new_n669), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n969), .B2(new_n328), .ZN(G1355gat));
endmodule


