

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739;

  XNOR2_X1 U368 ( .A(n391), .B(n348), .ZN(n390) );
  INV_X1 U369 ( .A(KEYINPUT35), .ZN(n348) );
  NAND2_X1 U370 ( .A1(n570), .A2(n656), .ZN(n552) );
  NOR2_X1 U371 ( .A1(n612), .A2(n445), .ZN(n449) );
  XNOR2_X1 U372 ( .A(n443), .B(n347), .ZN(n612) );
  XNOR2_X1 U373 ( .A(n717), .B(KEYINPUT4), .ZN(n347) );
  XNOR2_X1 U374 ( .A(n484), .B(n417), .ZN(n717) );
  XNOR2_X1 U375 ( .A(n418), .B(n434), .ZN(n484) );
  XNOR2_X1 U376 ( .A(G113), .B(KEYINPUT72), .ZN(n433) );
  NAND2_X1 U377 ( .A1(n620), .A2(G475), .ZN(n608) );
  NOR2_X2 U378 ( .A1(n687), .A2(n600), .ZN(n620) );
  INV_X1 U379 ( .A(n390), .ZN(n734) );
  NAND2_X1 U380 ( .A1(n390), .A2(n522), .ZN(n523) );
  NAND2_X1 U381 ( .A1(n405), .A2(n349), .ZN(n540) );
  NAND2_X1 U382 ( .A1(n524), .A2(n404), .ZN(n349) );
  NAND2_X2 U383 ( .A1(n563), .A2(n457), .ZN(n458) );
  INV_X1 U384 ( .A(n674), .ZN(n350) );
  XNOR2_X1 U385 ( .A(n496), .B(n495), .ZN(n674) );
  XNOR2_X1 U386 ( .A(n428), .B(n427), .ZN(n556) );
  XNOR2_X1 U387 ( .A(G119), .B(G116), .ZN(n436) );
  XNOR2_X1 U388 ( .A(KEYINPUT32), .B(n516), .ZN(n736) );
  BUF_X1 U389 ( .A(n667), .Z(n351) );
  NOR2_X1 U390 ( .A1(n528), .A2(n527), .ZN(n648) );
  XNOR2_X1 U391 ( .A(n386), .B(n387), .ZN(n671) );
  NOR2_X1 U392 ( .A1(n698), .A2(G902), .ZN(n428) );
  XNOR2_X1 U393 ( .A(n395), .B(n724), .ZN(n698) );
  XNOR2_X1 U394 ( .A(n442), .B(n356), .ZN(n395) );
  XNOR2_X1 U395 ( .A(n718), .B(KEYINPUT73), .ZN(n442) );
  XNOR2_X1 U396 ( .A(n422), .B(n421), .ZN(n718) );
  XNOR2_X1 U397 ( .A(n437), .B(G134), .ZN(n464) );
  XNOR2_X1 U398 ( .A(n435), .B(n436), .ZN(n418) );
  INV_X1 U399 ( .A(n433), .ZN(n435) );
  INV_X1 U400 ( .A(n423), .ZN(n437) );
  XNOR2_X1 U401 ( .A(G143), .B(G128), .ZN(n423) );
  INV_X2 U402 ( .A(G953), .ZN(n727) );
  XNOR2_X1 U403 ( .A(n556), .B(KEYINPUT1), .ZN(n667) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n487) );
  XOR2_X1 U405 ( .A(G137), .B(G140), .Z(n502) );
  XNOR2_X1 U406 ( .A(n389), .B(G125), .ZN(n467) );
  INV_X1 U407 ( .A(G146), .ZN(n389) );
  XNOR2_X1 U408 ( .A(n467), .B(n388), .ZN(n725) );
  INV_X1 U409 ( .A(KEYINPUT10), .ZN(n388) );
  OR2_X1 U410 ( .A1(n704), .A2(G902), .ZN(n387) );
  XNOR2_X1 U411 ( .A(n510), .B(n355), .ZN(n386) );
  NOR2_X1 U412 ( .A1(n637), .A2(n566), .ZN(n568) );
  NOR2_X1 U413 ( .A1(n662), .A2(n564), .ZN(n565) );
  NOR2_X1 U414 ( .A1(n580), .A2(n357), .ZN(n362) );
  AND2_X1 U415 ( .A1(n392), .A2(n390), .ZN(n375) );
  NOR2_X1 U416 ( .A1(n537), .A2(n538), .ZN(n374) );
  XNOR2_X1 U417 ( .A(n538), .B(KEYINPUT81), .ZN(n404) );
  XNOR2_X1 U418 ( .A(n424), .B(n464), .ZN(n486) );
  XOR2_X1 U419 ( .A(G137), .B(KEYINPUT5), .Z(n488) );
  NAND2_X1 U420 ( .A1(n385), .A2(n353), .ZN(n384) );
  XNOR2_X1 U421 ( .A(n583), .B(n369), .ZN(n385) );
  XOR2_X1 U422 ( .A(KEYINPUT102), .B(KEYINPUT104), .Z(n469) );
  XNOR2_X1 U423 ( .A(KEYINPUT103), .B(KEYINPUT101), .ZN(n468) );
  XNOR2_X1 U424 ( .A(G143), .B(G140), .ZN(n475) );
  XNOR2_X1 U425 ( .A(n381), .B(n467), .ZN(n380) );
  XNOR2_X1 U426 ( .A(n437), .B(n438), .ZN(n381) );
  XOR2_X1 U427 ( .A(KEYINPUT87), .B(KEYINPUT18), .Z(n440) );
  NOR2_X1 U428 ( .A1(n553), .A2(n670), .ZN(n558) );
  XOR2_X1 U429 ( .A(KEYINPUT85), .B(G107), .Z(n421) );
  INV_X1 U430 ( .A(G101), .ZN(n419) );
  XNOR2_X1 U431 ( .A(KEYINPUT16), .B(G122), .ZN(n417) );
  XNOR2_X1 U432 ( .A(n376), .B(n359), .ZN(n512) );
  NOR2_X1 U433 ( .A1(n531), .A2(n377), .ZN(n376) );
  NAND2_X1 U434 ( .A1(n414), .A2(KEYINPUT65), .ZN(n413) );
  INV_X1 U435 ( .A(n512), .ZN(n411) );
  NOR2_X1 U436 ( .A1(n351), .A2(n410), .ZN(n409) );
  NAND2_X1 U437 ( .A1(n350), .A2(n416), .ZN(n410) );
  INV_X1 U438 ( .A(KEYINPUT91), .ZN(n517) );
  XNOR2_X1 U439 ( .A(n506), .B(n505), .ZN(n704) );
  AND2_X1 U440 ( .A1(n569), .A2(n362), .ZN(n581) );
  INV_X1 U441 ( .A(KEYINPUT70), .ZN(n369) );
  XOR2_X1 U442 ( .A(G122), .B(G104), .Z(n474) );
  AND2_X1 U443 ( .A1(n589), .A2(n551), .ZN(n662) );
  XOR2_X1 U444 ( .A(KEYINPUT15), .B(G902), .Z(n445) );
  XNOR2_X1 U445 ( .A(G110), .B(G104), .ZN(n420) );
  XNOR2_X1 U446 ( .A(n486), .B(n394), .ZN(n724) );
  INV_X1 U447 ( .A(n502), .ZN(n394) );
  INV_X1 U448 ( .A(n445), .ZN(n600) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n452) );
  OR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n450) );
  NAND2_X1 U451 ( .A1(n482), .A2(n378), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U453 ( .A(KEYINPUT25), .ZN(n508) );
  NOR2_X1 U454 ( .A1(n670), .A2(n671), .ZN(n668) );
  XOR2_X1 U455 ( .A(G101), .B(G146), .Z(n491) );
  XNOR2_X1 U456 ( .A(n384), .B(n593), .ZN(n383) );
  INV_X1 U457 ( .A(n654), .ZN(n382) );
  XNOR2_X1 U458 ( .A(G128), .B(KEYINPUT93), .ZN(n499) );
  XNOR2_X1 U459 ( .A(G119), .B(G110), .ZN(n501) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n497) );
  INV_X1 U461 ( .A(KEYINPUT8), .ZN(n399) );
  NAND2_X1 U462 ( .A1(n727), .A2(G234), .ZN(n400) );
  XNOR2_X1 U463 ( .A(G116), .B(G107), .ZN(n459) );
  XNOR2_X1 U464 ( .A(n472), .B(n370), .ZN(n606) );
  XNOR2_X1 U465 ( .A(n442), .B(n379), .ZN(n443) );
  XNOR2_X1 U466 ( .A(n380), .B(n441), .ZN(n379) );
  NAND2_X1 U467 ( .A1(n354), .A2(n364), .ZN(n594) );
  NOR2_X1 U468 ( .A1(n589), .A2(n365), .ZN(n364) );
  INV_X1 U469 ( .A(n558), .ZN(n365) );
  NOR2_X1 U470 ( .A1(n562), .A2(n561), .ZN(n585) );
  INV_X1 U471 ( .A(n552), .ZN(n398) );
  AND2_X1 U472 ( .A1(n393), .A2(n407), .ZN(n366) );
  AND2_X1 U473 ( .A1(n554), .A2(n553), .ZN(n393) );
  NOR2_X1 U474 ( .A1(n512), .A2(n513), .ZN(n515) );
  XNOR2_X1 U475 ( .A(n532), .B(n371), .ZN(n649) );
  INV_X1 U476 ( .A(KEYINPUT31), .ZN(n371) );
  XNOR2_X1 U477 ( .A(n367), .B(KEYINPUT108), .ZN(n574) );
  NAND2_X1 U478 ( .A1(n412), .A2(n408), .ZN(n511) );
  NAND2_X1 U479 ( .A1(n411), .A2(n409), .ZN(n408) );
  AND2_X1 U480 ( .A1(n415), .A2(n413), .ZN(n412) );
  OR2_X1 U481 ( .A1(n674), .A2(n534), .ZN(n535) );
  NOR2_X1 U482 ( .A1(n526), .A2(n525), .ZN(n644) );
  XNOR2_X1 U483 ( .A(n703), .B(n704), .ZN(n368) );
  NOR2_X1 U484 ( .A1(n628), .A2(KEYINPUT44), .ZN(n352) );
  XOR2_X1 U485 ( .A(n592), .B(n591), .Z(n353) );
  NOR2_X1 U486 ( .A1(n571), .A2(n554), .ZN(n354) );
  XOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n355) );
  XOR2_X1 U488 ( .A(n426), .B(n425), .Z(n356) );
  AND2_X1 U489 ( .A1(n637), .A2(KEYINPUT47), .ZN(n357) );
  INV_X1 U490 ( .A(n392), .ZN(n628) );
  NAND2_X1 U491 ( .A1(n411), .A2(n366), .ZN(n392) );
  AND2_X1 U492 ( .A1(n655), .A2(n382), .ZN(n358) );
  XOR2_X1 U493 ( .A(n483), .B(KEYINPUT22), .Z(n359) );
  NAND2_X1 U494 ( .A1(n511), .A2(n671), .ZN(n635) );
  INV_X1 U495 ( .A(KEYINPUT65), .ZN(n416) );
  XOR2_X1 U496 ( .A(n700), .B(n699), .Z(n360) );
  XOR2_X1 U497 ( .A(KEYINPUT36), .B(KEYINPUT110), .Z(n361) );
  XOR2_X1 U498 ( .A(KEYINPUT84), .B(n604), .Z(n625) );
  AND2_X1 U499 ( .A1(n363), .A2(n625), .ZN(G54) );
  XNOR2_X1 U500 ( .A(n701), .B(n360), .ZN(n363) );
  XNOR2_X1 U501 ( .A(n479), .B(n471), .ZN(n370) );
  NAND2_X1 U502 ( .A1(n573), .A2(n572), .ZN(n367) );
  NOR2_X1 U503 ( .A1(n641), .A2(n577), .ZN(n579) );
  NOR2_X1 U504 ( .A1(n368), .A2(n705), .ZN(G66) );
  XNOR2_X1 U505 ( .A(n594), .B(KEYINPUT109), .ZN(n555) );
  NAND2_X1 U506 ( .A1(n374), .A2(n375), .ZN(n373) );
  NOR2_X1 U507 ( .A1(n649), .A2(n630), .ZN(n536) );
  NOR2_X1 U508 ( .A1(n554), .A2(n529), .ZN(n518) );
  NAND2_X1 U509 ( .A1(n373), .A2(n372), .ZN(n405) );
  NAND2_X1 U510 ( .A1(n352), .A2(n406), .ZN(n372) );
  INV_X1 U511 ( .A(n670), .ZN(n378) );
  NAND2_X1 U512 ( .A1(n383), .A2(n358), .ZN(n726) );
  NAND2_X1 U513 ( .A1(n521), .A2(n520), .ZN(n391) );
  NAND2_X1 U514 ( .A1(n396), .A2(n351), .ZN(n651) );
  XNOR2_X1 U515 ( .A(n397), .B(n361), .ZN(n396) );
  NAND2_X1 U516 ( .A1(n555), .A2(n398), .ZN(n397) );
  NOR2_X1 U517 ( .A1(n601), .A2(G902), .ZN(n466) );
  XNOR2_X1 U518 ( .A(n461), .B(n401), .ZN(n601) );
  XNOR2_X1 U519 ( .A(n402), .B(n463), .ZN(n401) );
  XNOR2_X1 U520 ( .A(n464), .B(n462), .ZN(n402) );
  INV_X1 U521 ( .A(n537), .ZN(n406) );
  INV_X1 U522 ( .A(n351), .ZN(n407) );
  OR2_X1 U523 ( .A1(n351), .A2(n674), .ZN(n414) );
  NAND2_X1 U524 ( .A1(n512), .A2(KEYINPUT65), .ZN(n415) );
  INV_X1 U525 ( .A(KEYINPUT76), .ZN(n567) );
  INV_X1 U526 ( .A(KEYINPUT78), .ZN(n578) );
  XNOR2_X1 U527 ( .A(n579), .B(n578), .ZN(n580) );
  INV_X1 U528 ( .A(n484), .ZN(n485) );
  XNOR2_X1 U529 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n593) );
  XNOR2_X1 U530 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U531 ( .A(n531), .B(n517), .ZN(n534) );
  XNOR2_X1 U532 ( .A(n622), .B(KEYINPUT111), .ZN(n623) );
  XNOR2_X1 U533 ( .A(n725), .B(n498), .ZN(n506) );
  XNOR2_X1 U534 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U535 ( .A(G131), .B(KEYINPUT4), .ZN(n424) );
  XOR2_X1 U536 ( .A(G146), .B(KEYINPUT92), .Z(n426) );
  NAND2_X1 U537 ( .A1(G227), .A2(n727), .ZN(n425) );
  XNOR2_X1 U538 ( .A(KEYINPUT71), .B(G469), .ZN(n427) );
  XOR2_X1 U539 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n430) );
  NAND2_X1 U540 ( .A1(G234), .A2(n600), .ZN(n429) );
  XNOR2_X1 U541 ( .A(n430), .B(n429), .ZN(n507) );
  NAND2_X1 U542 ( .A1(G221), .A2(n507), .ZN(n431) );
  XOR2_X1 U543 ( .A(KEYINPUT21), .B(n431), .Z(n432) );
  XNOR2_X1 U544 ( .A(KEYINPUT97), .B(n432), .ZN(n670) );
  XNOR2_X1 U545 ( .A(KEYINPUT86), .B(KEYINPUT3), .ZN(n434) );
  NAND2_X1 U546 ( .A1(G224), .A2(n727), .ZN(n438) );
  XNOR2_X1 U547 ( .A(KEYINPUT17), .B(KEYINPUT83), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U549 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n447) );
  NAND2_X1 U550 ( .A1(G210), .A2(n450), .ZN(n446) );
  XNOR2_X1 U551 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X2 U552 ( .A(n449), .B(n448), .ZN(n570) );
  NAND2_X1 U553 ( .A1(G214), .A2(n450), .ZN(n656) );
  XNOR2_X1 U554 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n451) );
  XNOR2_X2 U555 ( .A(n552), .B(n451), .ZN(n563) );
  XNOR2_X1 U556 ( .A(n452), .B(KEYINPUT14), .ZN(n454) );
  NAND2_X1 U557 ( .A1(G952), .A2(n454), .ZN(n453) );
  XOR2_X1 U558 ( .A(KEYINPUT90), .B(n453), .Z(n685) );
  NAND2_X1 U559 ( .A1(n727), .A2(n685), .ZN(n547) );
  NAND2_X1 U560 ( .A1(G902), .A2(n454), .ZN(n544) );
  INV_X1 U561 ( .A(n544), .ZN(n455) );
  NOR2_X1 U562 ( .A1(G898), .A2(n727), .ZN(n721) );
  NAND2_X1 U563 ( .A1(n455), .A2(n721), .ZN(n456) );
  NAND2_X1 U564 ( .A1(n547), .A2(n456), .ZN(n457) );
  XNOR2_X2 U565 ( .A(n458), .B(KEYINPUT0), .ZN(n531) );
  XOR2_X1 U566 ( .A(KEYINPUT7), .B(G122), .Z(n460) );
  XNOR2_X1 U567 ( .A(n460), .B(n459), .ZN(n463) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n462) );
  NAND2_X1 U569 ( .A1(G217), .A2(n497), .ZN(n461) );
  XNOR2_X1 U570 ( .A(KEYINPUT106), .B(G478), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n466), .B(n465), .ZN(n528) );
  XNOR2_X1 U572 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U573 ( .A(n725), .B(n470), .Z(n472) );
  NAND2_X1 U574 ( .A1(G214), .A2(n487), .ZN(n471) );
  XNOR2_X1 U575 ( .A(G113), .B(G131), .ZN(n473) );
  XNOR2_X1 U576 ( .A(n474), .B(n473), .ZN(n478) );
  XOR2_X1 U577 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n476) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U579 ( .A(n478), .B(n477), .Z(n479) );
  NOR2_X1 U580 ( .A1(G902), .A2(n606), .ZN(n481) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U582 ( .A(n481), .B(n480), .ZN(n527) );
  INV_X1 U583 ( .A(n527), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n528), .A2(n525), .ZN(n660) );
  INV_X1 U585 ( .A(n660), .ZN(n482) );
  XOR2_X1 U586 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n483) );
  XNOR2_X1 U587 ( .A(n486), .B(n485), .ZN(n494) );
  NAND2_X1 U588 ( .A1(n487), .A2(G210), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U590 ( .A(n490), .B(KEYINPUT99), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(n493), .ZN(n621) );
  NOR2_X1 U593 ( .A1(n621), .A2(G902), .ZN(n496) );
  INV_X1 U594 ( .A(G472), .ZN(n495) );
  NAND2_X1 U595 ( .A1(G221), .A2(n497), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n500) );
  XOR2_X1 U597 ( .A(n500), .B(n499), .Z(n504) );
  XNOR2_X1 U598 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U599 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U600 ( .A1(G217), .A2(n507), .ZN(n509) );
  XOR2_X1 U601 ( .A(KEYINPUT6), .B(n350), .Z(n554) );
  INV_X1 U602 ( .A(n554), .ZN(n513) );
  AND2_X1 U603 ( .A1(n671), .A2(n351), .ZN(n514) );
  NAND2_X1 U604 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U605 ( .A1(n635), .A2(n736), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n668), .A2(n667), .ZN(n529) );
  XNOR2_X1 U607 ( .A(KEYINPUT33), .B(n518), .ZN(n691) );
  NOR2_X1 U608 ( .A1(n534), .A2(n691), .ZN(n519) );
  XNOR2_X1 U609 ( .A(n519), .B(KEYINPUT34), .ZN(n521) );
  INV_X1 U610 ( .A(n528), .ZN(n526) );
  NAND2_X1 U611 ( .A1(n527), .A2(n526), .ZN(n575) );
  INV_X1 U612 ( .A(n575), .ZN(n520) );
  INV_X1 U613 ( .A(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U614 ( .A(n523), .B(KEYINPUT67), .ZN(n524) );
  INV_X1 U615 ( .A(n644), .ZN(n589) );
  XNOR2_X1 U616 ( .A(KEYINPUT107), .B(n648), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n350), .A2(n529), .ZN(n530) );
  XOR2_X1 U618 ( .A(KEYINPUT100), .B(n530), .Z(n678) );
  NOR2_X1 U619 ( .A1(n531), .A2(n678), .ZN(n532) );
  NAND2_X1 U620 ( .A1(n668), .A2(n556), .ZN(n533) );
  XNOR2_X1 U621 ( .A(n533), .B(KEYINPUT98), .ZN(n543) );
  NOR2_X1 U622 ( .A1(n543), .A2(n535), .ZN(n630) );
  NOR2_X1 U623 ( .A1(n662), .A2(n536), .ZN(n537) );
  INV_X1 U624 ( .A(KEYINPUT45), .ZN(n539) );
  XNOR2_X1 U625 ( .A(n540), .B(n539), .ZN(n711) );
  NAND2_X1 U626 ( .A1(n674), .A2(n656), .ZN(n541) );
  XNOR2_X1 U627 ( .A(KEYINPUT30), .B(n541), .ZN(n542) );
  NOR2_X1 U628 ( .A1(n543), .A2(n542), .ZN(n573) );
  NOR2_X1 U629 ( .A1(G900), .A2(n544), .ZN(n545) );
  NAND2_X1 U630 ( .A1(G953), .A2(n545), .ZN(n546) );
  NAND2_X1 U631 ( .A1(n547), .A2(n546), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n573), .A2(n557), .ZN(n549) );
  XOR2_X1 U633 ( .A(KEYINPUT38), .B(n570), .Z(n657) );
  INV_X1 U634 ( .A(n657), .ZN(n548) );
  NOR2_X1 U635 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U636 ( .A(n550), .B(KEYINPUT39), .ZN(n588) );
  NOR2_X1 U637 ( .A1(n588), .A2(n551), .ZN(n654) );
  INV_X1 U638 ( .A(n671), .ZN(n553) );
  INV_X1 U639 ( .A(n557), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n651), .B(KEYINPUT80), .ZN(n582) );
  INV_X1 U641 ( .A(n556), .ZN(n562) );
  NAND2_X1 U642 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U643 ( .A1(n350), .A2(n559), .ZN(n560) );
  XOR2_X1 U644 ( .A(KEYINPUT28), .B(n560), .Z(n561) );
  NAND2_X1 U645 ( .A1(n585), .A2(n563), .ZN(n637) );
  XNOR2_X1 U646 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n564) );
  XNOR2_X1 U647 ( .A(KEYINPUT77), .B(n565), .ZN(n566) );
  XNOR2_X1 U648 ( .A(n568), .B(n567), .ZN(n569) );
  INV_X1 U649 ( .A(n570), .ZN(n597) );
  NOR2_X1 U650 ( .A1(n571), .A2(n597), .ZN(n572) );
  NOR2_X2 U651 ( .A1(n575), .A2(n574), .ZN(n641) );
  NAND2_X1 U652 ( .A1(KEYINPUT47), .A2(n662), .ZN(n576) );
  XNOR2_X1 U653 ( .A(KEYINPUT79), .B(n576), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U655 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n592) );
  NAND2_X1 U656 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U657 ( .A1(n661), .A2(n660), .ZN(n584) );
  XNOR2_X1 U658 ( .A(KEYINPUT41), .B(n584), .ZN(n690) );
  INV_X1 U659 ( .A(n585), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n690), .A2(n586), .ZN(n587) );
  XNOR2_X1 U661 ( .A(n587), .B(KEYINPUT42), .ZN(n737) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT40), .ZN(n738) );
  NOR2_X1 U664 ( .A1(n737), .A2(n738), .ZN(n591) );
  NOR2_X1 U665 ( .A1(n351), .A2(n594), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n595), .A2(n656), .ZN(n596) );
  XNOR2_X1 U667 ( .A(KEYINPUT43), .B(n596), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n655) );
  NOR2_X1 U669 ( .A1(n711), .A2(n726), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT2), .ZN(n687) );
  BUF_X2 U671 ( .A(n620), .Z(n702) );
  NAND2_X1 U672 ( .A1(G478), .A2(n702), .ZN(n603) );
  INV_X1 U673 ( .A(n601), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n605) );
  NOR2_X1 U675 ( .A1(G952), .A2(n727), .ZN(n604) );
  INV_X1 U676 ( .A(n625), .ZN(n705) );
  AND2_X1 U677 ( .A1(n605), .A2(n625), .ZN(G63) );
  XNOR2_X1 U678 ( .A(n606), .B(KEYINPUT59), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n609), .A2(n625), .ZN(n611) );
  INV_X1 U681 ( .A(KEYINPUT60), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(G60) );
  NAND2_X1 U683 ( .A1(n620), .A2(G210), .ZN(n616) );
  XOR2_X1 U684 ( .A(n612), .B(KEYINPUT82), .Z(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n613) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n617), .A2(n625), .ZN(n619) );
  INV_X1 U688 ( .A(KEYINPUT56), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n619), .B(n618), .ZN(G51) );
  NAND2_X1 U690 ( .A1(n620), .A2(G472), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n621), .B(KEYINPUT62), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U694 ( .A(n627), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U695 ( .A(G101), .B(n628), .Z(G3) );
  NAND2_X1 U696 ( .A1(n630), .A2(n644), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(G104), .ZN(G6) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT26), .ZN(n634) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n632) );
  NAND2_X1 U700 ( .A1(n630), .A2(n648), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G9) );
  XOR2_X1 U703 ( .A(G110), .B(KEYINPUT113), .Z(n636) );
  XNOR2_X1 U704 ( .A(n635), .B(n636), .ZN(G12) );
  XOR2_X1 U705 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n639) );
  INV_X1 U706 ( .A(n637), .ZN(n642) );
  NAND2_X1 U707 ( .A1(n648), .A2(n642), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U709 ( .A(G128), .B(n640), .ZN(G30) );
  XOR2_X1 U710 ( .A(G143), .B(n641), .Z(G45) );
  NAND2_X1 U711 ( .A1(n642), .A2(n644), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(G146), .ZN(G48) );
  XOR2_X1 U713 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n646) );
  NAND2_X1 U714 ( .A1(n649), .A2(n644), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U716 ( .A(G113), .B(n647), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(G116), .ZN(G18) );
  XNOR2_X1 U719 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n652) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U721 ( .A(G125), .B(n653), .ZN(G27) );
  XOR2_X1 U722 ( .A(G134), .B(n654), .Z(G36) );
  XNOR2_X1 U723 ( .A(G140), .B(n655), .ZN(G42) );
  XOR2_X1 U724 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n697) );
  XOR2_X1 U725 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n684) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n658), .B(KEYINPUT118), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U731 ( .A(KEYINPUT119), .B(n665), .Z(n666) );
  NOR2_X1 U732 ( .A1(n691), .A2(n666), .ZN(n682) );
  NOR2_X1 U733 ( .A1(n668), .A2(n351), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT50), .B(n669), .Z(n676) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n672), .B(KEYINPUT49), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(KEYINPUT51), .B(n679), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n690), .A2(n680), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U743 ( .A(n684), .B(n683), .ZN(n686) );
  NAND2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n689) );
  BUF_X1 U745 ( .A(n687), .Z(n688) );
  NAND2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U748 ( .A(KEYINPUT121), .B(n692), .Z(n693) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n695), .A2(n727), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(G75) );
  XNOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT57), .ZN(n699) );
  NAND2_X1 U754 ( .A1(n702), .A2(G469), .ZN(n701) );
  NAND2_X1 U755 ( .A1(G217), .A2(n702), .ZN(n703) );
  NAND2_X1 U756 ( .A1(G224), .A2(KEYINPUT61), .ZN(n710) );
  INV_X1 U757 ( .A(G898), .ZN(n708) );
  AND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n706) );
  NOR2_X1 U759 ( .A1(KEYINPUT61), .A2(n706), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U762 ( .A1(G898), .A2(KEYINPUT61), .ZN(n712) );
  NAND2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n713), .A2(n727), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n716), .B(KEYINPUT125), .ZN(n723) );
  XNOR2_X1 U767 ( .A(n717), .B(n718), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n719), .B(KEYINPUT124), .ZN(n720) );
  NOR2_X1 U769 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U770 ( .A(n723), .B(n722), .Z(G69) );
  XNOR2_X1 U771 ( .A(n725), .B(n724), .ZN(n729) );
  XNOR2_X1 U772 ( .A(n726), .B(n729), .ZN(n728) );
  NAND2_X1 U773 ( .A1(n728), .A2(n727), .ZN(n733) );
  XNOR2_X1 U774 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U775 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U776 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U777 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U778 ( .A(G122), .B(KEYINPUT126), .ZN(n735) );
  XOR2_X1 U779 ( .A(n735), .B(n734), .Z(G24) );
  XNOR2_X1 U780 ( .A(G119), .B(n736), .ZN(G21) );
  XOR2_X1 U781 ( .A(G137), .B(n737), .Z(G39) );
  XNOR2_X1 U782 ( .A(G131), .B(KEYINPUT127), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n739), .B(n738), .ZN(G33) );
endmodule

