//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n541, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1087, new_n1088,
    new_n1089, new_n1090;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  OR2_X1    g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n452), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n459), .A3(G137), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  INV_X1    g046(.A(new_n459), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n472), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(new_n461), .B2(G114), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NOR2_X1   g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OR3_X1    g057(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n481), .B1(new_n480), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n465), .A2(new_n459), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n490), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n459), .A3(new_n492), .A4(new_n488), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n459), .A2(G126), .A3(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n485), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT71), .B1(new_n497), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(G88), .B1(G50), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT72), .ZN(G166));
  NAND3_X1  g088(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(G51), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(new_n505), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT73), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT7), .Z(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n510), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n508), .A2(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n516), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  NAND2_X1  g104(.A1(new_n508), .A2(G43), .ZN(new_n530));
  INV_X1    g105(.A(G81), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT74), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n510), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  XOR2_X1   g115(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n541));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G188));
  NAND3_X1  g119(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(KEYINPUT9), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n502), .A2(new_n503), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n506), .A2(G91), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n512), .B(new_n560), .ZN(G303));
  NAND3_X1  g136(.A1(new_n506), .A2(KEYINPUT77), .A3(G87), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n508), .A2(G49), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n516), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n562), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(G288));
  AND3_X1   g143(.A1(new_n504), .A2(G86), .A3(new_n505), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT78), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n554), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G651), .A3(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n506), .A2(G85), .B1(G47), .B2(new_n508), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n506), .A2(G92), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n507), .A2(KEYINPUT82), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n507), .A2(KEYINPUT82), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n590), .A2(G54), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n510), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G321));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G299), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G168), .B2(new_n598), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(G168), .B2(new_n598), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g182(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2100), .ZN(new_n611));
  AOI22_X1  g186(.A1(G123), .A2(new_n475), .B1(new_n473), .B2(G135), .ZN(new_n612));
  OAI221_X1 g187(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n615), .A2(G2096), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(G2096), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT84), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2438), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G1341), .B(G1348), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g209(.A(G2067), .B(G2678), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT18), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(KEYINPUT86), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT17), .Z(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n637), .B2(new_n636), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n635), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n638), .B1(new_n645), .B2(new_n637), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n641), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT87), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n648), .B(new_n650), .Z(G227));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT88), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT19), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  OR3_X1    g237(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT89), .B(G1981), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(G229));
  INV_X1    g246(.A(KEYINPUT105), .ZN(new_n672));
  NOR2_X1   g247(.A1(G16), .A2(G22), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(G166), .B2(G16), .ZN(new_n674));
  INV_X1    g249(.A(G1971), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(KEYINPUT91), .B1(G16), .B2(G23), .ZN(new_n677));
  OR3_X1    g252(.A1(KEYINPUT91), .A2(G16), .A3(G23), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n678), .C1(G288), .C2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT33), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(G6), .B(G305), .S(G16), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT90), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT32), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n676), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AOI22_X1  g264(.A1(G119), .A2(new_n475), .B1(new_n473), .B2(G131), .ZN(new_n690));
  OAI221_X1 g265(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n692), .S(G29), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT35), .B(G1991), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n679), .B1(new_n582), .B2(new_n584), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n679), .B2(G24), .ZN(new_n698));
  INV_X1    g273(.A(G1986), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(new_n698), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n689), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(KEYINPUT36), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n689), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT31), .B(G11), .ZN(new_n707));
  NAND2_X1  g282(.A1(G299), .A2(G16), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n679), .A2(KEYINPUT23), .A3(G20), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n710));
  INV_X1    g285(.A(G20), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT104), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT103), .B(G1956), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G27), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G164), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT30), .B(G28), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n717), .A2(G26), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n465), .A2(G116), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G104), .B2(G2105), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(G104), .A3(G2105), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n728), .A2(G2104), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n473), .A2(G140), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n475), .A2(G128), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G32), .ZN(new_n739));
  AOI22_X1  g314(.A1(G129), .A2(new_n475), .B1(new_n473), .B2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT26), .Z(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  AOI211_X1 g322(.A(new_n724), .B(new_n738), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AND4_X1   g323(.A1(new_n707), .A2(new_n716), .A3(new_n722), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G34), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n470), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT97), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  OR2_X1    g332(.A1(G29), .A2(G33), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n473), .A2(G139), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n760), .B(new_n761), .C1(new_n465), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(new_n717), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n757), .B(new_n767), .C1(new_n746), .C2(new_n747), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n615), .A2(new_n616), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n717), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n679), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n595), .B2(new_n679), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT92), .B(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n717), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n717), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT102), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n776), .B(new_n778), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n779), .A2(G2090), .B1(new_n720), .B2(new_n721), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n768), .A2(new_n770), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n754), .A2(new_n755), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(G2090), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n766), .B2(new_n765), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G171), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n749), .A2(new_n781), .A3(new_n782), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G21), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G168), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT98), .B(G1966), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n793), .B(new_n794), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n788), .A2(new_n785), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n706), .A2(new_n791), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n679), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n537), .B2(new_n679), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1341), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n672), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n796), .B(new_n790), .C1(new_n703), .C2(new_n705), .ZN(new_n803));
  INV_X1    g378(.A(new_n801), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n803), .A2(KEYINPUT105), .A3(new_n804), .A4(new_n795), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(G311));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n795), .ZN(G150));
  AOI22_X1  g382(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n510), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n508), .A2(G55), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n516), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n536), .B(new_n813), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n595), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n602), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n816), .B1(new_n822), .B2(G860), .ZN(G145));
  XNOR2_X1  g398(.A(new_n764), .B(new_n735), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n485), .A2(new_n494), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT106), .ZN(new_n826));
  AND3_X1   g401(.A1(new_n491), .A2(new_n826), .A3(new_n493), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n491), .B2(new_n493), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n744), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n824), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n475), .A2(G130), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT107), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n475), .A2(KEYINPUT107), .A3(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n473), .A2(G142), .ZN(new_n836));
  OAI221_X1 g411(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n465), .C2(G118), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n692), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT108), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n609), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n831), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n769), .B(new_n470), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n478), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(KEYINPUT110), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n831), .A2(new_n841), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(KEYINPUT110), .C2(new_n845), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT109), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n842), .B1(new_n849), .B2(new_n847), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n831), .A2(KEYINPUT109), .A3(new_n841), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g430(.A(G305), .B(KEYINPUT111), .ZN(new_n856));
  NAND2_X1  g431(.A1(G290), .A2(G166), .ZN(new_n857));
  NAND3_X1  g432(.A1(G303), .A2(new_n582), .A3(new_n584), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(G288), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(G288), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(new_n858), .ZN(new_n863));
  INV_X1    g438(.A(G288), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n856), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n859), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(KEYINPUT112), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT112), .B1(new_n862), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n595), .B(G299), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT41), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n817), .B(new_n604), .ZN(new_n875));
  MUX2_X1   g450(.A(new_n872), .B(new_n874), .S(new_n875), .Z(new_n876));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n877));
  INV_X1    g452(.A(new_n867), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n866), .B1(new_n865), .B2(new_n859), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n871), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n876), .B1(new_n871), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n814), .A2(new_n598), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n883), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n885), .ZN(G331));
  XNOR2_X1  g464(.A(G286), .B(G171), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n817), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(new_n872), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n873), .A2(new_n891), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n869), .A2(new_n870), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT112), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n878), .B2(new_n879), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n897), .A3(new_n868), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n898), .A3(new_n853), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n894), .A2(new_n898), .A3(new_n901), .A4(new_n853), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n900), .A2(new_n902), .B1(KEYINPUT114), .B2(KEYINPUT44), .ZN(new_n903));
  NOR2_X1   g478(.A1(KEYINPUT114), .A2(KEYINPUT44), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(G397));
  XOR2_X1   g480(.A(KEYINPUT115), .B(G1384), .Z(new_n906));
  AOI21_X1  g481(.A(KEYINPUT45), .B1(new_n829), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G40), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n466), .A2(new_n469), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n735), .B(new_n737), .ZN(new_n911));
  INV_X1    g486(.A(G1996), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n744), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT116), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n695), .A3(new_n691), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n916), .A2(new_n917), .B1(G2067), .B2(new_n735), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n919), .A2(new_n920), .A3(new_n910), .ZN(new_n921));
  INV_X1    g496(.A(new_n910), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT46), .B1(new_n922), .B2(new_n912), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT125), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(KEYINPUT46), .A3(new_n912), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n911), .A2(new_n745), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n924), .B(new_n926), .C1(new_n910), .C2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT47), .Z(new_n929));
  XNOR2_X1  g504(.A(new_n692), .B(new_n694), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n916), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(G290), .A2(G1986), .A3(new_n910), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT48), .Z(new_n933));
  AND2_X1   g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n921), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n829), .A2(KEYINPUT45), .A3(new_n906), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n466), .A2(new_n469), .A3(new_n908), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n495), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT117), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(G1971), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n829), .A2(new_n938), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n909), .B(new_n946), .C1(new_n947), .C2(KEYINPUT50), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(G2090), .ZN(new_n949));
  OAI21_X1  g524(.A(G8), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G8), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n942), .B(KEYINPUT117), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n675), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G2090), .B2(new_n948), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n951), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n958), .A3(G8), .ZN(new_n959));
  INV_X1    g534(.A(new_n574), .ZN(new_n960));
  OAI21_X1  g535(.A(G1981), .B1(new_n960), .B2(new_n569), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n962));
  OAI221_X1 g537(.A(new_n961), .B1(new_n962), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT49), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(G305), .A2(G1981), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(new_n962), .A3(KEYINPUT49), .A4(new_n961), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n829), .A2(new_n938), .A3(new_n909), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(G1976), .B2(new_n864), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n972), .B(new_n973), .C1(G1976), .C2(new_n864), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n953), .A2(new_n959), .A3(KEYINPUT63), .A4(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n948), .A2(G2084), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n909), .B1(new_n939), .B2(new_n940), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n947), .B2(new_n940), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n794), .ZN(new_n981));
  OAI21_X1  g556(.A(G8), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G286), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT63), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n976), .A2(G8), .A3(new_n956), .A4(new_n958), .ZN(new_n986));
  INV_X1    g561(.A(G1976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n971), .A2(new_n987), .A3(new_n864), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n985), .B(new_n986), .C1(new_n969), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n944), .A2(new_n721), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n992), .A2(new_n993), .B1(new_n785), .B2(new_n948), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n721), .A2(KEYINPUT53), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n980), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n991), .B(G301), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G286), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT122), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n982), .A2(KEYINPUT51), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n982), .A2(new_n999), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n978), .A2(new_n981), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n1002), .B2(new_n999), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n977), .A2(new_n983), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g580(.A(KEYINPUT62), .B(G301), .C1(new_n994), .C2(new_n996), .ZN(new_n1006));
  INV_X1    g581(.A(G1956), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n829), .B2(new_n938), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n495), .A2(new_n1008), .A3(new_n938), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n909), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1007), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n552), .A2(KEYINPUT57), .A3(new_n557), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n556), .A2(G651), .ZN(new_n1015));
  INV_X1    g590(.A(G91), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n516), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1017), .B2(new_n551), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n936), .A2(new_n941), .A3(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1012), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n968), .A2(G2067), .ZN(new_n1023));
  INV_X1    g598(.A(G1348), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n948), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1022), .A2(new_n820), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1019), .B1(new_n1012), .B2(new_n1021), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT61), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1012), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1032), .A2(KEYINPUT121), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1019), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n485), .A2(new_n494), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n491), .A2(new_n493), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT106), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n491), .A2(new_n826), .A3(new_n493), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT50), .B1(new_n1039), .B2(G1384), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1011), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1956), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n936), .A2(new_n941), .A3(new_n1020), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT121), .A3(new_n1032), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1031), .A2(new_n1033), .A3(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1046), .A2(KEYINPUT61), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1025), .A2(KEYINPUT60), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1025), .A2(KEYINPUT60), .A3(new_n820), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n820), .B1(new_n1025), .B2(KEYINPUT60), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1029), .B(new_n1030), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT58), .B(G1341), .Z(new_n1054));
  NAND2_X1  g629(.A1(new_n968), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n942), .B2(G1996), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1056), .B2(new_n537), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n537), .ZN(new_n1058));
  AND2_X1   g633(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1051), .A2(new_n1052), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1028), .B1(new_n1047), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n907), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(new_n936), .A3(new_n909), .A4(new_n995), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n994), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(G171), .B(KEYINPUT54), .Z(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n994), .A2(new_n996), .A3(new_n1066), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1006), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1005), .B1(new_n1071), .B2(new_n1004), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n959), .A2(new_n976), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n955), .B1(G2090), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n958), .B1(new_n1075), .B2(G8), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n990), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(G290), .B(new_n699), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n931), .B1(new_n910), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n935), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT127), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT127), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n935), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g660(.A1(new_n854), .A2(G319), .ZN(new_n1087));
  NOR2_X1   g661(.A1(new_n1087), .A2(G227), .ZN(new_n1088));
  NAND2_X1  g662(.A1(new_n900), .A2(new_n902), .ZN(new_n1089));
  INV_X1    g663(.A(G229), .ZN(new_n1090));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n633), .A4(new_n1090), .ZN(G225));
  INV_X1    g665(.A(G225), .ZN(G308));
endmodule


