//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT18), .A3(G131), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT18), .A2(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n191), .A2(new_n193), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n195), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n196), .A3(G125), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n200), .B2(new_n209), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n202), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n210), .C1(new_n200), .C2(new_n209), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n191), .B2(new_n193), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n191), .A2(new_n215), .A3(new_n193), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(KEYINPUT17), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n208), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G113), .B(G122), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n222), .A2(new_n223), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT88), .B1(new_n216), .B2(KEYINPUT17), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n214), .B(new_n220), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n228), .A3(new_n207), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(KEYINPUT89), .A3(new_n228), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n229), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(G475), .B1(new_n237), .B2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n217), .A2(new_n219), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n200), .B(KEYINPUT19), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n239), .B(new_n213), .C1(G146), .C2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n241), .A2(new_n207), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(new_n228), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n233), .A2(new_n234), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n233), .A2(new_n234), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n248));
  NOR2_X1   g062(.A1(G475), .A2(G902), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(KEYINPUT90), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n243), .B1(new_n236), .B2(new_n235), .ZN(new_n251));
  INV_X1    g065(.A(new_n249), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(new_n235), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n255), .B2(new_n244), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT90), .B1(new_n256), .B2(new_n248), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n238), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G902), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT93), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n190), .A2(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G134), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  INV_X1    g081(.A(G122), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G116), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT14), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT95), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT91), .B(G122), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n270), .B2(new_n269), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n267), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n269), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n267), .B(new_n278), .C1(new_n273), .C2(new_n274), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n266), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n262), .B1(new_n282), .B2(new_n263), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n263), .A2(new_n282), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT92), .ZN(new_n285));
  OAI21_X1  g099(.A(G134), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G107), .B1(new_n275), .B2(new_n269), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n279), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n262), .A2(new_n265), .A3(new_n263), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n290), .A2(KEYINPUT94), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(KEYINPUT94), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n281), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(G217), .A3(new_n188), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  AOI211_X1 g112(.A(new_n296), .B(new_n281), .C1(new_n291), .C2(new_n292), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n259), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G478), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G234), .ZN(new_n304));
  OAI211_X1 g118(.A(G952), .B(new_n188), .C1(new_n304), .C2(new_n187), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT96), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT21), .B(G898), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n259), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n292), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n290), .A2(KEYINPUT94), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n296), .B1(new_n314), .B2(new_n281), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n293), .A2(new_n297), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n302), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n259), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n303), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n258), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G469), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(new_n259), .ZN(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G140), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n188), .A2(G227), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT11), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n265), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n265), .A2(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n328), .A2(new_n330), .A3(new_n215), .A4(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n227), .A2(KEYINPUT76), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  AOI21_X1  g154(.A(G107), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT76), .B(G104), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n344), .B(KEYINPUT3), .C1(new_n345), .C2(G107), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n227), .A2(KEYINPUT3), .A3(G107), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n345), .B2(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n349), .A2(G101), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT78), .B(G101), .Z(new_n351));
  NAND4_X1  g165(.A1(new_n343), .A2(new_n351), .A3(new_n346), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n337), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(G101), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n202), .A2(G143), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n190), .A2(G146), .ZN(new_n359));
  AND2_X1   g173(.A1(KEYINPUT0), .A2(G128), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT64), .B1(new_n190), .B2(G146), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT0), .A2(G128), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n267), .A2(G104), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(G101), .C1(new_n341), .C2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n341), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT80), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n358), .A3(new_n359), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n358), .A2(new_n359), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n260), .B1(new_n358), .B2(KEYINPUT1), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND4_X1   g195(.A1(new_n352), .A2(new_n373), .A3(new_n375), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n352), .A2(new_n373), .A3(new_n375), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n190), .A2(G146), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n202), .B2(G143), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n377), .B1(new_n388), .B2(new_n380), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n377), .C1(new_n388), .C2(new_n380), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n392), .ZN(new_n393));
  OAI22_X1  g207(.A1(new_n382), .A2(KEYINPUT10), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n336), .B1(new_n370), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n368), .B1(new_n354), .B2(new_n356), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(new_n335), .A3(new_n394), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n326), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n370), .A2(new_n336), .A3(new_n395), .ZN(new_n400));
  INV_X1    g214(.A(new_n326), .ZN(new_n401));
  INV_X1    g215(.A(new_n373), .ZN(new_n402));
  INV_X1    g216(.A(new_n372), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n345), .B2(G107), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n371), .B1(new_n404), .B2(G101), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n389), .B1(new_n406), .B2(new_n352), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n335), .B1(new_n407), .B2(new_n382), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT12), .B1(new_n335), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI221_X1 g225(.A(new_n335), .B1(new_n409), .B2(KEYINPUT12), .C1(new_n407), .C2(new_n382), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n401), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(G902), .B1(new_n399), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n323), .B1(new_n415), .B2(new_n322), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n411), .A2(new_n412), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n398), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n400), .A2(KEYINPUT82), .A3(new_n413), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n326), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n398), .B2(new_n326), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n400), .A2(KEYINPUT83), .A3(new_n401), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n335), .B1(new_n397), .B2(new_n394), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(G469), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G221), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n295), .B2(new_n259), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n321), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT8), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n352), .A2(new_n373), .A3(new_n375), .ZN(new_n435));
  XNOR2_X1  g249(.A(G116), .B(G119), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n274), .A2(KEYINPUT5), .A3(G119), .ZN(new_n438));
  INV_X1    g252(.A(G113), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT2), .B(G113), .Z(new_n441));
  AOI22_X1  g255(.A1(new_n437), .A2(new_n440), .B1(new_n441), .B2(new_n436), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n435), .A2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n434), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n389), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n198), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n198), .B2(new_n367), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT85), .B(G224), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G953), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n448), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(new_n436), .ZN(new_n459));
  XOR2_X1   g273(.A(G116), .B(G119), .Z(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT2), .B(G113), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT65), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT65), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n355), .B2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n357), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n443), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n433), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n259), .B1(new_n458), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n433), .A2(KEYINPUT84), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n354), .B2(new_n356), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT6), .B(new_n475), .C1(new_n476), .C2(new_n443), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n443), .B1(new_n357), .B2(new_n468), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(new_n433), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n475), .B1(new_n476), .B2(new_n443), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n448), .B(new_n450), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT86), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n474), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  INV_X1    g305(.A(new_n477), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n471), .A2(KEYINPUT6), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(new_n481), .ZN(new_n494));
  INV_X1    g308(.A(new_n484), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n484), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n488), .A3(new_n474), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n490), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n432), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n265), .A2(G137), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n329), .A2(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n334), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n390), .A2(new_n392), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n367), .A2(new_n335), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n466), .B1(new_n510), .B2(KEYINPUT69), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT28), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT65), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n463), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n367), .A2(new_n335), .A3(KEYINPUT66), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT66), .B1(new_n367), .B2(new_n335), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n367), .A2(new_n335), .A3(KEYINPUT66), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n508), .A3(new_n517), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT28), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n515), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT29), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n192), .A2(G210), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT27), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n507), .A2(new_n389), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n509), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n466), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n525), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  INV_X1    g354(.A(new_n513), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n541), .A2(new_n542), .A3(new_n466), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n543), .B2(KEYINPUT28), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n530), .B(new_n535), .C1(KEYINPUT29), .C2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n523), .A2(new_n508), .A3(KEYINPUT30), .A4(new_n524), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n537), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n520), .A2(new_n547), .A3(KEYINPUT30), .A4(new_n508), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n526), .B1(new_n552), .B2(new_n466), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n534), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n545), .B(new_n259), .C1(KEYINPUT29), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n528), .B1(new_n525), .B2(new_n538), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n517), .A3(new_n513), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n528), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT70), .B1(new_n562), .B2(new_n535), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n564), .B(new_n534), .C1(new_n514), .C2(new_n559), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n552), .A2(new_n466), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n525), .A3(new_n535), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n553), .A2(new_n570), .A3(new_n535), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n558), .A2(new_n566), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n553), .B2(new_n535), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n517), .B1(new_n550), .B2(new_n551), .ZN(new_n574));
  NOR4_X1   g388(.A1(new_n574), .A2(KEYINPUT31), .A3(new_n526), .A4(new_n534), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n558), .B1(new_n576), .B2(new_n566), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n557), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n556), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n569), .A2(new_n571), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n564), .B1(new_n544), .B2(new_n534), .ZN(new_n582));
  INV_X1    g396(.A(new_n565), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT71), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n576), .A2(new_n558), .A3(new_n566), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT72), .B1(new_n587), .B2(new_n557), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n589));
  INV_X1    g403(.A(new_n557), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n589), .B(new_n590), .C1(new_n585), .C2(new_n586), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n580), .B1(new_n592), .B2(new_n579), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n212), .A2(new_n213), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n260), .A2(G119), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n260), .A2(G119), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT24), .B(G110), .Z(new_n599));
  INV_X1    g413(.A(KEYINPUT23), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n598), .A2(new_n599), .B1(new_n603), .B2(G110), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n598), .A2(new_n599), .B1(new_n603), .B2(G110), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n213), .A3(new_n203), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT22), .B(G137), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n429), .A2(new_n304), .A3(G953), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n605), .B2(new_n607), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n594), .B1(new_n616), .B2(G902), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT25), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n594), .B(KEYINPUT25), .C1(new_n616), .C2(G902), .ZN(new_n620));
  OAI21_X1  g434(.A(G217), .B1(new_n304), .B2(G902), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT73), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(G902), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT75), .B1(new_n593), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n578), .A2(new_n589), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n587), .A2(KEYINPUT72), .A3(new_n557), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n579), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n590), .B1(new_n585), .B2(new_n586), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n631), .A2(KEYINPUT32), .B1(G472), .B2(new_n555), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT75), .ZN(new_n634));
  INV_X1    g448(.A(new_n626), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n503), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n351), .ZN(G3));
  OAI21_X1  g452(.A(new_n259), .B1(new_n572), .B2(new_n577), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n430), .B(new_n626), .C1(new_n416), .C2(new_n427), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n592), .A2(KEYINPUT97), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n628), .A2(new_n640), .A3(new_n641), .A4(new_n629), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n488), .B1(new_n498), .B2(new_n474), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n489), .B(new_n473), .C1(new_n496), .C2(new_n497), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n501), .B(new_n311), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n317), .A2(KEYINPUT33), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n317), .A2(KEYINPUT33), .ZN(new_n650));
  OAI211_X1 g464(.A(G478), .B(new_n259), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(KEYINPUT98), .A2(G478), .ZN(new_n652));
  AND2_X1   g466(.A1(KEYINPUT98), .A2(G478), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n300), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n258), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n642), .A2(new_n645), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G6));
  NAND2_X1  g475(.A1(new_n303), .A2(new_n319), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n251), .A2(KEYINPUT20), .A3(new_n252), .ZN(new_n663));
  INV_X1    g477(.A(new_n253), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n662), .B(new_n238), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n648), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n642), .A2(new_n645), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n608), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n624), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n623), .A2(new_n672), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n628), .A2(new_n640), .A3(new_n629), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n502), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  OAI21_X1  g491(.A(new_n501), .B1(new_n646), .B2(new_n647), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n309), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n306), .B1(G900), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT100), .Z(new_n682));
  NOR2_X1   g496(.A1(new_n665), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n430), .B1(new_n416), .B2(new_n427), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n673), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n633), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n678), .B1(new_n630), .B2(new_n632), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n685), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(G128), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G30));
  NOR2_X1   g507(.A1(new_n646), .A2(new_n647), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n258), .A2(new_n662), .ZN(new_n697));
  INV_X1    g511(.A(new_n501), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n697), .A2(new_n698), .A3(new_n673), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n682), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n699), .B1(new_n701), .B2(KEYINPUT40), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(KEYINPUT40), .B2(new_n701), .ZN(new_n703));
  INV_X1    g517(.A(G472), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n553), .A2(new_n534), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(G902), .B1(new_n527), .B2(new_n534), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI221_X1 g522(.A(new_n630), .B1(new_n579), .B2(new_n578), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT103), .B(G143), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G45));
  INV_X1    g526(.A(new_n682), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n655), .A2(new_n258), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n688), .A2(new_n684), .A3(new_n673), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT104), .B(G146), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G48));
  INV_X1    g532(.A(new_n414), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n401), .B1(new_n400), .B2(new_n425), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n259), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n322), .B(new_n259), .C1(new_n719), .C2(new_n720), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n430), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n657), .A2(new_n633), .A3(new_n635), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n666), .A2(new_n633), .A3(new_n635), .A4(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  INV_X1    g544(.A(new_n725), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n678), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n633), .A2(new_n732), .A3(new_n321), .A4(new_n673), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  XNOR2_X1  g548(.A(new_n557), .B(KEYINPUT105), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n529), .A2(new_n534), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n581), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n585), .B2(new_n586), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n635), .B(new_n737), .C1(new_n738), .C2(new_n704), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n725), .A2(new_n311), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n698), .B(new_n697), .C1(new_n490), .C2(new_n499), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  OAI211_X1 g558(.A(new_n673), .B(new_n737), .C1(new_n738), .C2(new_n704), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n714), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND2_X1  g562(.A1(new_n578), .A2(new_n579), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n626), .B1(new_n632), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n490), .A2(new_n501), .A3(new_n499), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n421), .A2(G469), .A3(new_n426), .ZN(new_n753));
  INV_X1    g567(.A(new_n323), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n723), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n416), .A2(KEYINPUT106), .A3(new_n427), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n431), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n750), .A2(new_n759), .A3(KEYINPUT42), .A4(new_n715), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n633), .A2(new_n635), .A3(new_n759), .A4(new_n715), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n763), .B1(new_n761), .B2(KEYINPUT107), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n760), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT108), .B(G131), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G33));
  NAND4_X1  g581(.A1(new_n633), .A2(new_n635), .A3(new_n759), .A4(new_n683), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT109), .B(G134), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G36));
  NAND2_X1  g584(.A1(new_n421), .A2(new_n426), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n322), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n754), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n778), .B1(new_n322), .B2(new_n415), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n430), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n258), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n655), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n783), .B2(KEYINPUT111), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n655), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n784), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n592), .A2(new_n640), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n673), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n751), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n781), .A2(new_n795), .A3(new_n700), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NOR4_X1   g612(.A1(new_n633), .A2(new_n635), .A3(new_n714), .A4(new_n751), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  AOI211_X1 g615(.A(new_n801), .B(new_n430), .C1(new_n779), .C2(new_n780), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  OR2_X1    g618(.A1(new_n724), .A2(KEYINPUT49), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n724), .A2(KEYINPUT49), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n626), .A2(new_n698), .A3(new_n430), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OR4_X1    g622(.A1(new_n709), .A2(new_n696), .A3(new_n787), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n751), .A2(new_n731), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT119), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n791), .A2(new_n307), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n750), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT48), .ZN(new_n815));
  INV_X1    g629(.A(new_n739), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n732), .ZN(new_n818));
  OAI211_X1 g632(.A(G952), .B(new_n188), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n656), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n709), .A2(new_n306), .A3(new_n626), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n811), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n695), .A2(new_n698), .A3(new_n725), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT50), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n822), .A2(new_n782), .A3(new_n654), .A4(new_n651), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n813), .A2(new_n640), .A3(new_n673), .A4(new_n737), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n800), .A2(new_n802), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n431), .B2(new_n724), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n817), .A2(new_n751), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT118), .Z(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n824), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n835), .A2(KEYINPUT120), .A3(KEYINPUT51), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT120), .B1(new_n835), .B2(KEYINPUT51), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n689), .A2(new_n633), .A3(new_n679), .A4(new_n685), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n689), .B1(new_n688), .B2(new_n685), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n716), .B(new_n747), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n758), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n673), .A2(new_n682), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n709), .A2(new_n742), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT52), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n747), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n687), .B2(new_n690), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n847), .A3(new_n852), .A4(new_n716), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n238), .B(new_n713), .C1(new_n664), .C2(new_n663), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n662), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n303), .A2(KEYINPUT113), .A3(new_n319), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n684), .A3(new_n673), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n751), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n633), .A2(new_n862), .B1(new_n759), .B2(new_n746), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n768), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(KEYINPUT114), .A3(new_n768), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n502), .A2(new_n674), .B1(new_n741), .B2(new_n742), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n658), .A2(new_n869), .A3(new_n733), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n637), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n648), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n782), .A2(new_n859), .A3(new_n858), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n642), .A2(new_n645), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n726), .A3(new_n729), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n868), .A2(new_n765), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n691), .A2(new_n747), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n855), .A2(new_n879), .A3(KEYINPUT53), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n854), .B2(new_n878), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n854), .A2(new_n878), .A3(new_n884), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n878), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n849), .A2(new_n853), .A3(new_n881), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n637), .A2(new_n876), .A3(new_n870), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT115), .A3(new_n765), .A4(new_n868), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n887), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI211_X1 g708(.A(KEYINPUT116), .B(new_n886), .C1(new_n894), .C2(new_n883), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n884), .ZN(new_n896));
  INV_X1    g710(.A(new_n887), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT54), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n841), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n809), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NAND2_X1  g717(.A1(new_n882), .A2(new_n885), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G902), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(G210), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT56), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n483), .B(new_n495), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n188), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n911), .A2(new_n916), .ZN(G51));
  NAND2_X1  g731(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n886), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n323), .B(KEYINPUT57), .ZN(new_n920));
  AOI22_X1  g734(.A1(new_n919), .A2(new_n920), .B1(new_n399), .B2(new_n414), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n905), .A2(new_n776), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n921), .B2(KEYINPUT122), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n926), .A2(KEYINPUT123), .A3(new_n251), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n926), .B2(new_n251), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n912), .B1(new_n926), .B2(new_n251), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n895), .A2(new_n900), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n649), .A2(new_n650), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n919), .B(new_n932), .C1(new_n649), .C2(new_n650), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n913), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n904), .A2(new_n671), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n904), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n913), .B(new_n943), .C1(new_n944), .C2(new_n615), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT61), .Z(G66));
  NOR2_X1   g760(.A1(new_n449), .A2(new_n308), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n188), .ZN(new_n948));
  INV_X1    g762(.A(new_n891), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n188), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n494), .B1(G898), .B2(new_n188), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(G69));
  XOR2_X1   g766(.A(new_n552), .B(new_n240), .Z(new_n953));
  INV_X1    g767(.A(new_n844), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n710), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n627), .A2(new_n636), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n701), .B(new_n751), .C1(new_n656), .C2(new_n873), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n797), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n956), .A2(new_n803), .A3(new_n957), .A4(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n953), .B1(new_n962), .B2(new_n188), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n750), .A2(new_n742), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n781), .A2(new_n700), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n965), .A2(new_n768), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n966), .A2(new_n803), .A3(new_n765), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n797), .A2(new_n954), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n797), .A2(new_n970), .A3(new_n954), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n967), .A2(new_n972), .A3(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n188), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n953), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n963), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n977), .B2(new_n979), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  AOI221_X4 g799(.A(new_n963), .B1(new_n981), .B2(new_n985), .C1(new_n977), .C2(new_n979), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G72));
  NAND3_X1  g801(.A1(new_n975), .A2(new_n891), .A3(new_n976), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  AOI21_X1  g804(.A(new_n554), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n990), .B1(new_n962), .B2(new_n949), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n912), .B1(new_n992), .B2(new_n705), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n706), .A2(new_n554), .A3(new_n990), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(new_n894), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n991), .A2(new_n995), .ZN(G57));
endmodule


