//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT1), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n217), .A2(new_n219), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n219), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(KEYINPUT25), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n215), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n223), .A2(new_n224), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n222), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n214), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n243), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n212), .B1(new_n236), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G227gat), .ZN(new_n250));
  INV_X1    g049(.A(G233gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n221), .A2(new_n219), .A3(new_n222), .ZN(new_n254));
  AND2_X1   g053(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n214), .A2(new_n213), .B1(new_n255), .B2(G190gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n224), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n235), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n220), .B2(KEYINPUT23), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(new_n219), .A3(new_n226), .A4(new_n227), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n212), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n243), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT28), .B1(new_n242), .B2(new_n243), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n214), .B(new_n240), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n253), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT34), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n271));
  NOR3_X1   g070(.A1(new_n236), .A2(new_n248), .A3(new_n212), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n263), .B1(new_n262), .B2(new_n266), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n252), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n249), .A2(new_n267), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n252), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT69), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G15gat), .ZN(new_n282));
  INV_X1    g081(.A(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n270), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n276), .B2(new_n278), .ZN(new_n288));
  INV_X1    g087(.A(new_n271), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT67), .B1(new_n277), .B2(new_n252), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n275), .B(new_n253), .C1(new_n249), .C2(new_n267), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n268), .B(KEYINPUT34), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n284), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n286), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n288), .B1(new_n286), .B2(new_n294), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n298));
  INV_X1    g097(.A(G141gat), .ZN(new_n299));
  INV_X1    g098(.A(G148gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n305));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G155gat), .B(G162gat), .Z(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  XNOR2_X1  g109(.A(G155gat), .B(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT2), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n311), .A2(new_n301), .A3(new_n314), .A4(new_n306), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G197gat), .ZN(new_n319));
  INV_X1    g118(.A(G204gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  NOR2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT70), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  INV_X1    g129(.A(G218gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(new_n324), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n322), .ZN(new_n336));
  OAI22_X1  g135(.A1(new_n335), .A2(new_n336), .B1(new_n326), .B2(KEYINPUT22), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT70), .B1(new_n326), .B2(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n332), .A2(new_n329), .A3(new_n324), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n318), .A2(new_n341), .A3(KEYINPUT80), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT80), .B1(new_n318), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n334), .A2(new_n340), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT3), .B1(new_n345), .B2(new_n317), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n309), .A2(new_n315), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(G228gat), .B(G233gat), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n298), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n318), .A2(new_n341), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n318), .A2(new_n341), .A3(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n310), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(new_n347), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G22gat), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n362));
  INV_X1    g161(.A(new_n334), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n363), .B2(KEYINPUT79), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT3), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n309), .A2(new_n367), .A3(new_n315), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n351), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n356), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n360), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n361), .B1(new_n360), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT82), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n344), .A2(new_n349), .A3(new_n298), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT81), .B1(new_n355), .B2(new_n358), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G22gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n361), .A3(new_n371), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT31), .B(G50gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n297), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT87), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n262), .A2(new_n266), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n262), .A2(new_n396), .A3(new_n266), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n317), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n230), .A2(new_n235), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n246), .A2(new_n247), .ZN(new_n402));
  INV_X1    g201(.A(new_n241), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n401), .A2(new_n257), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT72), .B1(new_n404), .B2(new_n399), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT72), .ZN(new_n406));
  INV_X1    g205(.A(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n345), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n397), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n407), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n407), .A2(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n341), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n393), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n399), .B1(new_n395), .B2(new_n397), .ZN(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n345), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n405), .A2(new_n408), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n399), .B2(new_n398), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n392), .C1(new_n421), .C2(new_n345), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n410), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n419), .A4(new_n392), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n204), .A2(KEYINPUT74), .A3(new_n211), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT74), .B1(new_n204), .B2(new_n211), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n428), .B(new_n316), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n212), .A2(new_n347), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT78), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n366), .A2(new_n263), .A3(new_n435), .A4(new_n368), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(KEYINPUT4), .C1(new_n212), .C2(new_n347), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n347), .B1(new_n429), .B2(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(new_n434), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n432), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(new_n441), .ZN(new_n447));
  INV_X1    g246(.A(new_n432), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n212), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n204), .A2(new_n211), .A3(KEYINPUT74), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n348), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n452), .B2(new_n434), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n366), .A2(new_n263), .A3(KEYINPUT4), .A4(new_n368), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n435), .B1(new_n212), .B2(new_n347), .ZN(new_n457));
  AND4_X1   g256(.A1(new_n456), .A2(new_n431), .A3(new_n432), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT77), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(new_n458), .C1(new_n447), .C2(new_n454), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n442), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT0), .ZN(new_n465));
  XNOR2_X1  g264(.A(G57gat), .B(G85gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  INV_X1    g268(.A(new_n467), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n470), .B(new_n442), .C1(new_n460), .C2(new_n462), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n467), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n427), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n297), .A2(new_n386), .A3(new_n475), .A4(new_n387), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n389), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n388), .A2(KEYINPUT35), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n473), .ZN(new_n482));
  INV_X1    g281(.A(new_n427), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n386), .B2(new_n387), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n386), .A2(new_n485), .A3(new_n387), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n297), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n440), .A2(new_n431), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n448), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n452), .A2(new_n448), .A3(new_n434), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n432), .B1(new_n440), .B2(new_n431), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n467), .B1(new_n499), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT40), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n463), .B2(new_n467), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(new_n496), .A3(new_n448), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n470), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n499), .A2(new_n496), .A3(new_n495), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT84), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n498), .A2(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n504), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n427), .A2(new_n503), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT85), .ZN(new_n515));
  INV_X1    g314(.A(new_n422), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n412), .A2(new_n341), .A3(new_n414), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT86), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n421), .A2(new_n345), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n517), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT38), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n416), .B1(new_n519), .B2(new_n392), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n393), .A2(KEYINPUT37), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n416), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n519), .B1(new_n424), .B2(new_n419), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT38), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n525), .A2(new_n472), .A3(new_n473), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n386), .A2(new_n387), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n489), .B(new_n492), .C1(new_n515), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n481), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n536), .A2(KEYINPUT89), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n539), .A2(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G43gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n283), .A2(G50gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT15), .ZN(new_n546));
  INV_X1    g345(.A(G29gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n536), .ZN(new_n550));
  NOR3_X1   g349(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n549), .A2(KEYINPUT15), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n542), .A2(new_n546), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G99gat), .B(G106gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT7), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(G85gat), .A3(G92gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n556), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n565), .A3(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI221_X1 g368(.A(KEYINPUT17), .B1(new_n548), .B2(new_n552), .C1(new_n542), .C2(new_n546), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n573));
  INV_X1    g372(.A(new_n568), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n566), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n553), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI211_X1 g377(.A(KEYINPUT98), .B(new_n573), .C1(new_n553), .C2(new_n575), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n572), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n581), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n586), .B(new_n571), .C1(new_n578), .C2(new_n579), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n582), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT94), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G57gat), .B(G64gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n593), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n596), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G57gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(G64gat), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G57gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(KEYINPUT95), .A3(G64gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n361), .A2(G15gat), .ZN(new_n618));
  INV_X1    g417(.A(G15gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(G22gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT90), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G1gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(G1gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G15gat), .B(G22gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT16), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(G8gat), .ZN(new_n630));
  INV_X1    g429(.A(G8gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n622), .A2(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n625), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n614), .B2(new_n613), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n617), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G183gat), .B(G211gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT97), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n636), .B(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n590), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n556), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n602), .A2(new_n612), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n575), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n602), .A2(new_n612), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n569), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n575), .A2(KEYINPUT10), .A3(new_n612), .A4(new_n602), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n575), .B(new_n651), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(new_n656), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  INV_X1    g463(.A(new_n662), .ZN(new_n665));
  INV_X1    g464(.A(new_n656), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n653), .B2(new_n654), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n658), .A2(new_n656), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT100), .B(new_n665), .C1(new_n667), .C2(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT18), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n634), .A2(new_n555), .A3(new_n570), .ZN(new_n674));
  NAND2_X1  g473(.A1(G229gat), .A2(G233gat), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT91), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n553), .B(new_n676), .C1(new_n630), .C2(new_n633), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n629), .A2(G8gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n632), .A2(new_n631), .A3(new_n625), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n676), .B1(new_n681), .B2(new_n553), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n674), .B(new_n675), .C1(new_n678), .C2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT92), .B1(new_n681), .B2(new_n553), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT92), .ZN(new_n685));
  INV_X1    g484(.A(new_n553), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n634), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n684), .B(new_n687), .C1(new_n678), .C2(new_n682), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n675), .B(KEYINPUT13), .Z(new_n689));
  AOI22_X1  g488(.A1(new_n673), .A2(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n553), .B1(new_n630), .B2(new_n633), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT91), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n677), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(KEYINPUT18), .A3(new_n675), .A4(new_n674), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT93), .B1(new_n683), .B2(new_n673), .ZN(new_n695));
  XNOR2_X1  g494(.A(G113gat), .B(G141gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT88), .B(G197gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT11), .B(G169gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT12), .Z(new_n701));
  OAI211_X1 g500(.A(new_n690), .B(new_n694), .C1(new_n695), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n673), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT93), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n689), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n706), .A3(new_n694), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n645), .A2(new_n672), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n535), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n482), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n623), .ZN(G1324gat));
  INV_X1    g512(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n427), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT16), .B(G8gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT101), .ZN(new_n719));
  MUX2_X1   g518(.A(KEYINPUT102), .B(new_n717), .S(new_n719), .Z(new_n720));
  NOR2_X1   g519(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n716), .B1(new_n715), .B2(G8gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n714), .A2(new_n427), .A3(new_n719), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(G1325gat));
  INV_X1    g523(.A(new_n297), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n711), .A2(G15gat), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n714), .A2(new_n491), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(G15gat), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT103), .ZN(G1326gat));
  AND3_X1   g528(.A1(new_n386), .A2(new_n485), .A3(new_n387), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n486), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  INV_X1    g534(.A(new_n590), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n481), .B2(new_n534), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n702), .A2(new_n708), .ZN(new_n738));
  INV_X1    g537(.A(new_n644), .ZN(new_n739));
  INV_X1    g538(.A(new_n672), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n482), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n547), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n491), .B1(new_n731), .B2(new_n484), .ZN(new_n748));
  INV_X1    g547(.A(new_n442), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n446), .A2(new_n443), .A3(new_n441), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT76), .B1(new_n453), .B2(KEYINPUT5), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n459), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n461), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n455), .A2(KEYINPUT77), .A3(new_n459), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n501), .B1(new_n755), .B2(new_n470), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n511), .B1(new_n510), .B2(new_n504), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT84), .B(KEYINPUT40), .C1(new_n498), .C2(new_n500), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT85), .B1(new_n760), .B2(new_n427), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT85), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n514), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n532), .B(new_n530), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n478), .A2(new_n480), .B1(new_n748), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n747), .B1(new_n765), .B2(new_n736), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n535), .A2(KEYINPUT44), .A3(new_n590), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n741), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT104), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n766), .A2(new_n767), .A3(new_n770), .A4(new_n741), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(new_n744), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n746), .B1(new_n772), .B2(new_n547), .ZN(G1328gat));
  NOR3_X1   g572(.A1(new_n742), .A2(G36gat), .A3(new_n483), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT46), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n769), .A2(new_n427), .A3(new_n771), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n538), .ZN(G1329gat));
  OAI21_X1  g576(.A(G43gat), .B1(new_n768), .B2(new_n492), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n742), .A2(G43gat), .A3(new_n725), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n769), .A2(new_n491), .A3(new_n771), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(G43gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g583(.A(G50gat), .B1(new_n768), .B2(new_n532), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n742), .A2(G50gat), .A3(new_n732), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(KEYINPUT48), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n731), .A3(new_n771), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(G50gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g590(.A1(new_n535), .A2(new_n645), .A3(new_n740), .A4(new_n738), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n482), .B(KEYINPUT105), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(new_n605), .ZN(G1332gat));
  NOR2_X1   g594(.A1(new_n483), .A2(new_n672), .ZN(new_n796));
  AND4_X1   g595(.A1(new_n535), .A2(new_n645), .A3(new_n738), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  AND2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(G1333gat));
  OR3_X1    g600(.A1(new_n792), .A2(KEYINPUT106), .A3(new_n725), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT106), .B1(new_n792), .B2(new_n725), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n594), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n792), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(G71gat), .A3(new_n491), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT50), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1334gat));
  NOR2_X1   g610(.A1(new_n792), .A2(new_n732), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(new_n595), .ZN(G1335gat));
  NOR2_X1   g612(.A1(new_n709), .A2(new_n739), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n766), .A2(new_n767), .A3(new_n740), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815), .B2(new_n482), .ZN(new_n816));
  AND4_X1   g615(.A1(KEYINPUT51), .A2(new_n535), .A3(new_n590), .A4(new_n814), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n737), .B2(new_n814), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n744), .A2(new_n563), .A3(new_n740), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1336gat));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(KEYINPUT107), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n796), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n564), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n564), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n766), .A2(new_n767), .A3(new_n814), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(KEYINPUT107), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n824), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n535), .A2(new_n590), .A3(new_n814), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n814), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(G92gat), .B1(new_n837), .B2(new_n796), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n830), .A3(new_n823), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n832), .A2(new_n839), .ZN(G1337gat));
  OAI21_X1  g639(.A(G99gat), .B1(new_n815), .B2(new_n492), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n725), .A2(G99gat), .A3(new_n672), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n819), .B2(new_n842), .ZN(G1338gat));
  NOR3_X1   g642(.A1(new_n532), .A2(G106gat), .A3(new_n672), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT109), .Z(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n817), .B2(new_n818), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT110), .ZN(new_n847));
  XNOR2_X1  g646(.A(KEYINPUT108), .B(G106gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n815), .B2(new_n732), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n837), .A2(new_n850), .A3(new_n845), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT53), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n837), .B2(new_n844), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n815), .B2(new_n532), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(G1339gat));
  NAND3_X1  g656(.A1(new_n645), .A2(new_n738), .A3(new_n672), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n700), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n688), .A2(new_n689), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n675), .B1(new_n693), .B2(new_n674), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n703), .A2(new_n706), .A3(new_n701), .A4(new_n694), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT113), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n653), .A2(new_n666), .A3(new_n654), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT112), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n653), .A2(new_n873), .A3(new_n666), .A4(new_n654), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n872), .A2(new_n657), .A3(KEYINPUT54), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n662), .B1(new_n667), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT55), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(KEYINPUT55), .A3(new_n877), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n590), .A2(new_n663), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n870), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT114), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n881), .A2(new_n663), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n709), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n672), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n736), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n881), .A2(new_n663), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT55), .B1(new_n875), .B2(new_n877), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n590), .A3(new_n869), .A4(new_n867), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n884), .A2(new_n890), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n860), .B1(new_n897), .B2(new_n644), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n731), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n744), .A2(new_n483), .A3(new_n297), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(G113gat), .B1(new_n903), .B2(new_n738), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n898), .A2(new_n793), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n389), .A2(new_n476), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n427), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n709), .A2(new_n207), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT115), .Z(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n904), .A2(new_n911), .ZN(G1340gat));
  AOI21_X1  g711(.A(G120gat), .B1(new_n908), .B2(new_n740), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n672), .A2(new_n209), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n902), .B2(new_n914), .ZN(G1341gat));
  OAI21_X1  g714(.A(G127gat), .B1(new_n903), .B2(new_n644), .ZN(new_n916));
  INV_X1    g715(.A(G127gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n908), .A2(new_n917), .A3(new_n739), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1342gat));
  OR4_X1    g718(.A1(G134gat), .A2(new_n907), .A3(new_n427), .A4(new_n736), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n921));
  OAI21_X1  g720(.A(G134gat), .B1(new_n903), .B2(new_n736), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1343gat));
  NOR2_X1   g723(.A1(new_n491), .A2(new_n532), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n427), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n299), .A3(new_n709), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n897), .A2(new_n644), .ZN(new_n929));
  INV_X1    g728(.A(new_n860), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT57), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n531), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT57), .B1(new_n898), .B2(new_n732), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n491), .A2(new_n482), .A3(new_n427), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G141gat), .B1(new_n936), .B2(new_n738), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(G1344gat));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n941), .B(G148gat), .C1(new_n936), .C2(new_n672), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n590), .B1(new_n886), .B2(new_n888), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n883), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n887), .B1(new_n893), .B2(new_n709), .ZN(new_n946));
  OAI211_X1 g745(.A(KEYINPUT118), .B(new_n894), .C1(new_n946), .C2(new_n590), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(new_n644), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n858), .B(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n732), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT119), .B1(new_n952), .B2(KEYINPUT57), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n894), .B1(new_n946), .B2(new_n590), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n739), .B1(new_n955), .B2(new_n943), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n950), .B1(new_n956), .B2(new_n947), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n954), .B(new_n932), .C1(new_n957), .C2(new_n732), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n931), .A2(KEYINPUT57), .A3(new_n531), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n935), .A2(new_n740), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n300), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n942), .B1(new_n962), .B2(new_n941), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n927), .A2(new_n300), .A3(new_n740), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1345gat));
  NAND3_X1  g764(.A1(new_n927), .A2(new_n312), .A3(new_n739), .ZN(new_n966));
  OAI21_X1  g765(.A(G155gat), .B1(new_n936), .B2(new_n644), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1346gat));
  OAI21_X1  g767(.A(G162gat), .B1(new_n936), .B2(new_n736), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n483), .A2(new_n313), .A3(new_n590), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n926), .B2(new_n970), .ZN(G1347gat));
  NAND2_X1  g770(.A1(new_n793), .A2(new_n427), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(new_n725), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n973), .A2(new_n899), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(G169gat), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n975), .A2(new_n976), .A3(new_n738), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n931), .A2(KEYINPUT120), .A3(new_n482), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT120), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n898), .B2(new_n744), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(new_n427), .A3(new_n906), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n709), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n977), .B1(new_n983), .B2(new_n976), .ZN(G1348gat));
  INV_X1    g783(.A(G176gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n982), .A2(new_n985), .A3(new_n740), .ZN(new_n986));
  OAI21_X1  g785(.A(G176gat), .B1(new_n975), .B2(new_n672), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1349gat));
  NAND3_X1  g787(.A1(new_n982), .A2(new_n242), .A3(new_n739), .ZN(new_n989));
  OAI21_X1  g788(.A(G183gat), .B1(new_n975), .B2(new_n644), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g790(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n991), .B(new_n992), .ZN(G1350gat));
  AOI21_X1  g792(.A(new_n243), .B1(new_n974), .B2(new_n590), .ZN(new_n994));
  XNOR2_X1  g793(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n982), .A2(new_n243), .A3(new_n590), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n997), .A2(KEYINPUT122), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n997), .A2(KEYINPUT122), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(G1351gat));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n427), .A3(new_n925), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(KEYINPUT124), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n981), .A2(new_n1003), .A3(new_n427), .A4(new_n925), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n1002), .A2(new_n319), .A3(new_n709), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT125), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n972), .A2(new_n491), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n960), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(G197gat), .B1(new_n1008), .B2(new_n738), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1006), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1352gat));
  AND4_X1   g811(.A1(new_n320), .A2(new_n981), .A3(new_n796), .A4(new_n925), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g814(.A(G204gat), .B1(new_n1008), .B2(new_n672), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(G1353gat));
  NAND4_X1  g817(.A1(new_n1002), .A2(new_n330), .A3(new_n739), .A4(new_n1004), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1020));
  NAND4_X1  g819(.A1(new_n960), .A2(new_n1020), .A3(new_n739), .A4(new_n1007), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1021), .A2(G211gat), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n960), .A2(new_n739), .A3(new_n1007), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(KEYINPUT126), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AND4_X1   g824(.A1(KEYINPUT63), .A2(new_n1024), .A3(G211gat), .A4(new_n1021), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(G1354gat));
  NOR3_X1   g826(.A1(new_n1008), .A2(new_n331), .A3(new_n736), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1002), .A2(new_n590), .A3(new_n1004), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1029), .A2(new_n331), .ZN(new_n1030));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1029), .A2(KEYINPUT127), .A3(new_n331), .ZN(new_n1033));
  AOI21_X1  g832(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(G1355gat));
endmodule


