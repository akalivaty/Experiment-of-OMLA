//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  OR2_X1    g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G43gat), .A2(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(KEYINPUT91), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT91), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n207), .A3(new_n204), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n203), .A2(KEYINPUT92), .A3(new_n202), .A4(new_n204), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT14), .B(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n205), .B2(KEYINPUT15), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n217), .A2(new_n220), .B1(new_n206), .B2(new_n208), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT93), .B(KEYINPUT17), .Z(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n209), .A2(new_n210), .B1(new_n214), .B2(new_n216), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT17), .B1(new_n226), .B2(new_n221), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G1gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G1gat), .B2(new_n228), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n225), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n226), .A2(new_n221), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n231), .B(G8gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G141gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G197gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT11), .B(G169gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n238), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n233), .B1(new_n226), .B2(new_n221), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n238), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(new_n235), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n241), .A2(new_n246), .A3(new_n247), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n239), .A2(new_n240), .B1(new_n249), .B2(new_n252), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n246), .B1(new_n256), .B2(new_n247), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n262), .A2(new_n264), .B1(G183gat), .B2(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT27), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT27), .B(G183gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G190gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  AOI21_X1  g079(.A(G190gat), .B1(new_n267), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT28), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n265), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT64), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(G183gat), .A3(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AND4_X1   g098(.A1(KEYINPUT25), .A2(new_n296), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n290), .A2(new_n303), .A3(new_n291), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n301), .A2(KEYINPUT65), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT65), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n283), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT1), .ZN(new_n311));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT25), .A4(new_n299), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n292), .B2(new_n289), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n284), .A2(new_n288), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n319), .B(new_n320), .C1(G183gat), .C2(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT25), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n315), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n301), .A2(KEYINPUT65), .A3(new_n306), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n313), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n283), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n314), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT34), .Z(new_n332));
  XNOR2_X1  g131(.A(G15gat), .B(G43gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT71), .ZN(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(new_n328), .B2(new_n330), .ZN(new_n340));
  AOI211_X1 g139(.A(KEYINPUT69), .B(new_n329), .C1(new_n314), .C2(new_n327), .ZN(new_n341));
  OAI211_X1 g140(.A(KEYINPUT32), .B(new_n338), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n332), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n273), .A2(new_n280), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n267), .A2(new_n280), .ZN(new_n347));
  INV_X1    g146(.A(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n275), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n277), .ZN(new_n351));
  AOI221_X4 g150(.A(new_n313), .B1(new_n351), .B2(new_n265), .C1(new_n323), .C2(new_n324), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n326), .B1(new_n325), .B2(new_n283), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n330), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT69), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n339), .A3(new_n330), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n336), .B1(new_n357), .B2(new_n337), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT70), .B1(new_n357), .B2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n360), .B(new_n361), .C1(new_n355), .C2(new_n356), .ZN(new_n362));
  OAI211_X1 g161(.A(KEYINPUT72), .B(new_n358), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT32), .B1(new_n340), .B2(new_n341), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n360), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT72), .B1(new_n368), .B2(new_n358), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n345), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n358), .B1(new_n359), .B2(new_n362), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n363), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT74), .B1(new_n376), .B2(new_n345), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n259), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n371), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(KEYINPUT74), .A3(new_n345), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT75), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n344), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n378), .A2(new_n381), .B1(new_n332), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n309), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT77), .Z(new_n388));
  NAND3_X1  g187(.A1(new_n325), .A2(KEYINPUT78), .A3(new_n283), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n283), .B1(new_n322), .B2(new_n317), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n387), .B1(new_n392), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(G197gat), .ZN(new_n397));
  INV_X1    g196(.A(G204gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n401), .B(new_n402), .ZN(new_n404));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405));
  MUX2_X1   g204(.A(new_n403), .B(new_n404), .S(new_n405), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n387), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n409), .A3(new_n389), .ZN(new_n410));
  INV_X1    g209(.A(new_n388), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT30), .B1(new_n419), .B2(KEYINPUT80), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n424));
  INV_X1    g223(.A(new_n417), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(KEYINPUT79), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n420), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434));
  OR2_X1    g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(G141gat), .B(G148gat), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n434), .B(new_n435), .C1(new_n436), .C2(KEYINPUT2), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  INV_X1    g237(.A(G148gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G141gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT82), .B(G141gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n434), .B1(new_n435), .B2(KEYINPUT2), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n437), .A2(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n437), .A2(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n406), .A2(new_n409), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n449), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n406), .B1(new_n452), .B2(new_n409), .ZN(new_n453));
  OR3_X1    g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n451), .B1(new_n450), .B2(new_n453), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n455), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n451), .B(new_n458), .C1(new_n450), .C2(new_n453), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n433), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n433), .A3(new_n459), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G22gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n460), .A3(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n446), .B(new_n326), .ZN(new_n475));
  NAND2_X1  g274(.A1(G225gat), .A2(G233gat), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n477));
  NOR3_X1   g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n446), .A2(new_n313), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT4), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n326), .B1(new_n446), .B2(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n452), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n476), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n477), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n488), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n478), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT0), .ZN(new_n493));
  XNOR2_X1  g292(.A(G57gat), .B(G85gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n493), .B(new_n494), .Z(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n495), .B(KEYINPUT88), .Z(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n491), .B2(new_n496), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n473), .A2(new_n474), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n384), .A2(new_n429), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n379), .A2(new_n380), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n383), .A2(new_n332), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n473), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n491), .A2(new_n496), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n497), .B1(new_n509), .B2(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n429), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT35), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n466), .A2(new_n461), .A3(new_n467), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n460), .B1(new_n470), .B2(new_n465), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n468), .A2(KEYINPUT87), .A3(new_n471), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n484), .A2(new_n485), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n475), .A2(new_n476), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT39), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n498), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n524), .B(new_n525), .C1(KEYINPUT39), .C2(new_n522), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n499), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT89), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n472), .B1(new_n428), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n424), .A2(KEYINPUT37), .A3(new_n426), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n417), .B1(new_n414), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT38), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n539));
  INV_X1    g338(.A(new_n406), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n535), .B1(new_n395), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n412), .A2(new_n540), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT38), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n503), .A2(new_n544), .A3(new_n419), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n538), .A2(KEYINPUT90), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n533), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n379), .A2(KEYINPUT75), .A3(new_n380), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT75), .B1(new_n379), .B2(new_n380), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n507), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n506), .A2(new_n507), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT36), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n521), .A2(new_n548), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n258), .B1(new_n513), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(G71gat), .ZN(new_n558));
  INV_X1    g357(.A(G78gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n562), .ZN(new_n567));
  OR2_X1    g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n564), .A3(new_n560), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  INV_X1    g372(.A(G231gat), .ZN(new_n574));
  INV_X1    g373(.A(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n573), .A2(new_n577), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n579), .A2(new_n580), .A3(G127gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n237), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(G127gat), .B1(new_n579), .B2(new_n580), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G127gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n580), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n583), .B1(new_n589), .B2(new_n581), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  INV_X1    g390(.A(G155gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT96), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n586), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n586), .B2(new_n590), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT97), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT98), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT7), .B1(new_n607), .B2(new_n605), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n608), .B(new_n612), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n609), .ZN(new_n621));
  INV_X1    g420(.A(new_n609), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT100), .B1(new_n622), .B2(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n617), .A2(new_n624), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n225), .A2(new_n227), .A3(new_n628), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n236), .A2(new_n627), .B1(KEYINPUT41), .B2(new_n599), .ZN(new_n630));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n604), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n631), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n603), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n597), .A2(new_n598), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT102), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n563), .A2(new_n565), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n564), .B1(new_n570), .B2(new_n560), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n625), .B2(new_n626), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n617), .A2(new_n624), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n617), .A2(new_n624), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n572), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n651), .A3(KEYINPUT101), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n627), .A2(new_n653), .A3(new_n572), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n644), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n643), .A3(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n641), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n556), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n510), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT103), .B(G1gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  NOR2_X1   g472(.A1(new_n670), .A2(new_n429), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n232), .B2(new_n674), .ZN(new_n677));
  MUX2_X1   g476(.A(new_n676), .B(new_n677), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n552), .A2(new_n679), .A3(new_n554), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n552), .B2(new_n554), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n670), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n384), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n670), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n519), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n513), .A2(new_n555), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n640), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n635), .A2(new_n639), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n513), .B2(new_n555), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n597), .A2(new_n598), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(new_n258), .A3(new_n667), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n510), .ZN(new_n701));
  INV_X1    g500(.A(new_n510), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n695), .A2(new_n215), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n700), .B2(new_n429), .ZN(new_n706));
  INV_X1    g505(.A(new_n698), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n668), .A3(new_n640), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n429), .A2(G36gat), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n556), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n552), .A2(new_n554), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n693), .A2(new_n713), .A3(new_n699), .A4(new_n696), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n708), .A2(G43gat), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n556), .A2(new_n384), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n680), .A2(new_n681), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n693), .A2(new_n720), .A3(new_n699), .A4(new_n696), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n717), .B1(new_n721), .B2(G43gat), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n715), .A2(new_n719), .B1(new_n722), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n693), .A2(new_n472), .A3(new_n699), .A4(new_n696), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G50gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n519), .A2(G50gat), .A3(new_n708), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n556), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n693), .A2(new_n520), .A3(new_n699), .A4(new_n696), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n729), .A2(G50gat), .B1(new_n556), .B2(new_n726), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g530(.A(new_n258), .ZN(new_n732));
  NOR4_X1   g531(.A1(new_n732), .A2(new_n707), .A3(new_n668), .A4(new_n640), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n690), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n690), .A2(KEYINPUT105), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n702), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n738), .A2(new_n429), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n738), .B2(new_n682), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n736), .A2(new_n558), .A3(new_n384), .A4(new_n737), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n519), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n559), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n732), .A2(new_n698), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n667), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n697), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n510), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(KEYINPUT108), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(KEYINPUT108), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n695), .B(new_n757), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n691), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n764), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n610), .A3(new_n702), .A4(new_n667), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n761), .A2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n429), .A2(G92gat), .A3(new_n668), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n693), .A2(new_n428), .A3(new_n696), .A4(new_n759), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n768), .A2(new_n771), .B1(new_n773), .B2(G92gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n760), .B2(new_n682), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n668), .A2(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n768), .A2(new_n384), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n473), .A2(G106gat), .A3(new_n668), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n693), .A2(new_n472), .A3(new_n696), .A4(new_n759), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n693), .A2(new_n520), .A3(new_n696), .A4(new_n759), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n768), .A2(new_n784), .B1(new_n790), .B2(G106gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n791), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n644), .C1(new_n655), .C2(new_n657), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n664), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n655), .A2(new_n644), .A3(new_n657), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT54), .B(new_n658), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT55), .B(new_n796), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n235), .B1(new_n234), .B2(new_n238), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n248), .A2(new_n238), .A3(new_n251), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n245), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n245), .C1(new_n805), .C2(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n254), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n694), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n803), .A2(new_n666), .A3(new_n804), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(KEYINPUT112), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n804), .A2(new_n666), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n640), .A2(new_n254), .A3(new_n808), .A4(new_n810), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n801), .B2(new_n802), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n732), .A3(new_n666), .A4(new_n804), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n668), .A2(new_n811), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n694), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n698), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n641), .A2(new_n258), .A3(new_n668), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT109), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n641), .A2(KEYINPUT109), .A3(new_n668), .A4(new_n258), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n793), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n813), .A2(KEYINPUT112), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n818), .A3(new_n815), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n640), .B1(new_n821), .B2(new_n823), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n707), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n520), .B1(new_n833), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n428), .A2(new_n510), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n384), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(G113gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(new_n258), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n510), .B1(new_n833), .B2(new_n839), .ZN(new_n845));
  INV_X1    g644(.A(new_n508), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n428), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n732), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(new_n843), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n842), .A2(new_n851), .A3(new_n668), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n667), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n851), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n587), .A3(new_n698), .ZN(new_n855));
  OAI21_X1  g654(.A(G127gat), .B1(new_n842), .B2(new_n707), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NAND2_X1  g656(.A1(new_n429), .A2(new_n640), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n847), .A2(G134gat), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n842), .B2(new_n694), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NAND3_X1  g663(.A1(new_n552), .A2(new_n554), .A3(new_n841), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n552), .A2(new_n867), .A3(new_n554), .A4(new_n841), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n520), .B(KEYINPUT57), .C1(new_n826), .C2(new_n832), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n473), .B1(new_n833), .B2(new_n839), .ZN(new_n871));
  XNOR2_X1  g670(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n441), .B1(new_n875), .B2(new_n258), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n472), .B(new_n845), .C1(new_n680), .C2(new_n681), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n428), .ZN(new_n878));
  INV_X1    g677(.A(G141gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n732), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n881), .B(new_n882), .ZN(G1344gat));
  NOR2_X1   g682(.A1(new_n439), .A2(KEYINPUT59), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n875), .B2(new_n668), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n887));
  AOI21_X1  g686(.A(new_n258), .B1(new_n801), .B2(new_n802), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n822), .B1(new_n816), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n834), .B(new_n835), .C1(new_n889), .C2(new_n640), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n793), .B(new_n832), .C1(new_n890), .C2(new_n707), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT113), .B1(new_n838), .B2(new_n831), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n472), .B(new_n873), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(new_n827), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n825), .A2(new_n813), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n707), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(new_n519), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(new_n667), .A3(new_n866), .A4(new_n868), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT118), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G148gat), .B1(new_n900), .B2(KEYINPUT118), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n886), .B(new_n887), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n869), .A2(new_n906), .A3(new_n667), .A4(new_n899), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(G148gat), .A3(new_n901), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n886), .B1(new_n908), .B2(new_n887), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n885), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n878), .A2(new_n439), .A3(new_n667), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(G155gat), .B1(new_n875), .B2(new_n707), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n878), .A2(new_n592), .A3(new_n698), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n875), .B2(new_n694), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n858), .A2(G162gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n877), .B2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n508), .A2(new_n429), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n920), .B(new_n510), .C1(new_n892), .C2(new_n891), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n732), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n429), .A2(new_n702), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n384), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n925), .A2(KEYINPUT121), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(KEYINPUT121), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n840), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n294), .A3(new_n258), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n923), .A2(new_n929), .ZN(G1348gat));
  OAI21_X1  g729(.A(G176gat), .B1(new_n928), .B2(new_n668), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n667), .A2(new_n295), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n921), .B2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n928), .B2(new_n707), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n698), .A2(new_n272), .A3(new_n274), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n921), .C2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n348), .A3(new_n640), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n928), .A2(new_n694), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n348), .B1(new_n941), .B2(KEYINPUT61), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n940), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n939), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  OAI21_X1  g745(.A(new_n924), .B1(new_n680), .B2(new_n681), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n871), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n732), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n896), .A2(new_n707), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n827), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT57), .B1(new_n953), .B2(new_n520), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n871), .B2(new_n873), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n947), .B2(KEYINPUT124), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n957), .B(new_n924), .C1(new_n680), .C2(new_n681), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n258), .A2(new_n397), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n956), .A2(new_n667), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n398), .B1(new_n962), .B2(KEYINPUT126), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(KEYINPUT126), .B2(new_n962), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n949), .A2(G204gat), .A3(new_n668), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(KEYINPUT125), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n964), .B(new_n967), .C1(new_n965), .C2(new_n968), .ZN(G1353gat));
  OR3_X1    g768(.A1(new_n949), .A2(G211gat), .A3(new_n707), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n956), .A2(KEYINPUT127), .A3(new_n698), .A4(new_n958), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(G211gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n973), .A2(new_n698), .A3(new_n899), .A4(new_n958), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  AND4_X1   g776(.A1(KEYINPUT63), .A2(new_n976), .A3(G211gat), .A4(new_n971), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n950), .A2(new_n980), .A3(new_n640), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n959), .A2(new_n640), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n980), .ZN(G1355gat));
endmodule


