//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND2_X1  g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n470), .A2(G137), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n469), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n469), .A2(new_n471), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n470), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n471), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n467), .B2(new_n468), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n489), .B(new_n494), .C1(new_n468), .C2(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n512), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(new_n510), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(new_n522), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(new_n510), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n523), .A2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n512), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n521), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n523), .A2(G52), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n512), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n521), .A2(G81), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT75), .B(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n523), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT77), .ZN(G188));
  AOI22_X1  g130(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n512), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(G91), .B2(new_n521), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n523), .A2(new_n559), .A3(G53), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n518), .A2(G543), .A3(new_n519), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(G299));
  NAND4_X1  g142(.A1(new_n518), .A2(G49), .A3(G543), .A4(new_n519), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n520), .C2(new_n570), .ZN(G288));
  NAND4_X1  g146(.A1(new_n518), .A2(G86), .A3(new_n510), .A4(new_n519), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n515), .A2(new_n517), .B1(KEYINPUT6), .B2(new_n512), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n574), .A2(new_n575), .A3(G86), .A4(new_n510), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n508), .B2(new_n509), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n518), .A2(G48), .A3(G543), .A4(new_n519), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n577), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n521), .A2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n512), .C2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n574), .A2(G92), .A3(new_n510), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n510), .A2(G66), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n512), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G54), .B2(new_n523), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G286), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g177(.A(G299), .B(KEYINPUT80), .Z(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n471), .A2(G2104), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n476), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G2100), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT81), .ZN(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(G111), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G2105), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n480), .A2(G123), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  AOI211_X1 g200(.A(new_n623), .B(new_n625), .C1(G135), .C2(new_n470), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n620), .A2(new_n626), .B1(new_n617), .B2(G2100), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n619), .B(new_n627), .C1(new_n620), .C2(new_n626), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n647), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n648), .ZN(new_n654));
  INV_X1    g229(.A(new_n647), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n648), .B(new_n656), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n651), .B(new_n654), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n646), .A2(new_n655), .A3(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n650), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT20), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n664), .A2(new_n666), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n669), .A3(new_n667), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n674), .C1(new_n669), .C2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G11), .ZN(new_n682));
  INV_X1    g257(.A(G28), .ZN(new_n683));
  AOI21_X1  g258(.A(G29), .B1(new_n683), .B2(KEYINPUT30), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(KEYINPUT30), .B2(new_n683), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n688), .B1(new_n626), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NOR2_X1   g269(.A1(G164), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G27), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G2078), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G2072), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n689), .A2(G33), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT93), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n470), .A2(G139), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n704), .C1(new_n471), .C2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G29), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n693), .B(new_n698), .C1(new_n699), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n694), .A2(G26), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n470), .A2(G140), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n480), .A2(G128), .ZN(new_n713));
  OR2_X1    g288(.A1(G104), .A2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n689), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2067), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n708), .B(new_n719), .C1(new_n699), .C2(new_n707), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n689), .A2(G32), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n613), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n480), .A2(G129), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  AND3_X1   g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(new_n689), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT27), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1996), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G34), .ZN(new_n730));
  AOI22_X1  g305(.A1(G160), .A2(G29), .B1(new_n694), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G2084), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G2084), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n697), .B2(new_n696), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n548), .B2(new_n735), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n732), .B(new_n734), .C1(G1341), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n720), .A2(new_n729), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT98), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT23), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G1956), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G4), .A2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT91), .Z(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n597), .B2(new_n735), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(G1348), .Z(new_n749));
  NOR2_X1   g324(.A1(new_n737), .A2(G1341), .ZN(new_n750));
  NAND2_X1  g325(.A1(G168), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G16), .B2(G21), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT95), .B(G1966), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT94), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n750), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n752), .B2(new_n754), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n739), .A2(new_n745), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G24), .B(G290), .S(G16), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT89), .B(G1986), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n470), .A2(G131), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n480), .A2(G119), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n765));
  OAI221_X1 g340(.A(G2104), .B1(G107), .B2(new_n471), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n761), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G25), .B(new_n767), .S(new_n692), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT35), .B(G1991), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G6), .B(G305), .S(G16), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n735), .A2(G22), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G166), .B2(new_n735), .ZN(new_n775));
  INV_X1    g350(.A(G1971), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n735), .A2(G23), .ZN(new_n778));
  INV_X1    g353(.A(G288), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n735), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n773), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n760), .B(new_n770), .C1(new_n783), .C2(KEYINPUT34), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(KEYINPUT34), .B2(new_n783), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(KEYINPUT36), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n786), .A2(KEYINPUT36), .ZN(new_n789));
  OR3_X1    g364(.A1(new_n785), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n692), .A2(G35), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n692), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2090), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n735), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n735), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT97), .ZN(new_n797));
  INV_X1    g372(.A(G1961), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n757), .A2(new_n788), .A3(new_n790), .A4(new_n800), .ZN(G150));
  INV_X1    g376(.A(G150), .ZN(G311));
  NOR2_X1   g377(.A1(new_n597), .A2(new_n606), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT38), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(new_n512), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n521), .A2(G93), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n523), .A2(G55), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n547), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n547), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n804), .B(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(KEYINPUT39), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(KEYINPUT39), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n814), .A2(new_n815), .A3(G860), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(G860), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT99), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  OR2_X1    g394(.A1(new_n816), .A2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n504), .A2(KEYINPUT101), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n499), .A2(new_n822), .A3(new_n503), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n471), .A2(G138), .ZN(new_n824));
  OR2_X1    g399(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n825));
  NAND2_X1  g400(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT72), .B(KEYINPUT4), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n497), .B(KEYINPUT100), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT100), .B1(new_n496), .B2(new_n497), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n821), .B(new_n823), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n717), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n726), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n726), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n480), .A2(G130), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n471), .A2(G118), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G142), .B2(new_n470), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n615), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n767), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n839), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(new_n478), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n626), .ZN(new_n849));
  AOI21_X1  g424(.A(G37), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n847), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g427(.A1(G299), .A2(new_n598), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n597), .B(new_n558), .C1(new_n565), .C2(new_n566), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(G299), .A2(KEYINPUT103), .A3(new_n598), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n856), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n859), .A3(new_n855), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n857), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n608), .B(new_n812), .ZN(new_n863));
  MUX2_X1   g438(.A(new_n861), .B(new_n862), .S(new_n863), .Z(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT42), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT42), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(G288), .B(KEYINPUT104), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(G290), .B(G303), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n869), .B(new_n870), .Z(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(KEYINPUT105), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n873), .A3(new_n866), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(G868), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT106), .B1(new_n809), .B2(new_n601), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n875), .B2(new_n878), .ZN(G295));
  AOI21_X1  g454(.A(new_n877), .B1(new_n875), .B2(new_n878), .ZN(G331));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n810), .A2(new_n811), .A3(G301), .ZN(new_n882));
  AOI21_X1  g457(.A(G301), .B1(new_n810), .B2(new_n811), .ZN(new_n883));
  OAI21_X1  g458(.A(G286), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n812), .A2(G171), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n810), .A2(new_n811), .A3(G301), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(G168), .A3(new_n886), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n884), .A2(new_n887), .B1(new_n856), .B2(new_n857), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n861), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n858), .B2(new_n860), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT107), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n895), .A3(new_n871), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n871), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n894), .B2(new_n888), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n881), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n889), .A2(new_n859), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n853), .A2(new_n855), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n862), .B1(new_n889), .B2(new_n859), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n909), .A2(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT44), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n902), .B2(new_n903), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n881), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n918), .ZN(G397));
  INV_X1    g494(.A(KEYINPUT63), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n832), .A2(KEYINPUT45), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G40), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n478), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(G1384), .B1(new_n498), .B2(new_n505), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n922), .A2(KEYINPUT110), .A3(new_n924), .A4(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n776), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n832), .A2(KEYINPUT111), .A3(new_n921), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n832), .B2(new_n921), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G2090), .ZN(new_n937));
  NAND2_X1  g512(.A1(G160), .A2(G40), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT116), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n925), .A2(KEYINPUT116), .A3(new_n939), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n936), .A2(new_n937), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G8), .ZN(new_n946));
  NAND2_X1  g521(.A1(G303), .A2(G8), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n821), .A2(new_n823), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n498), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n954), .B2(new_n829), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n955), .B2(G1384), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n832), .A2(KEYINPUT111), .A3(new_n921), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n939), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n926), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n925), .B2(new_n939), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n938), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n937), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n950), .B1(new_n933), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n948), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n957), .A3(new_n924), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n779), .A2(G1976), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT114), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n967), .A2(G8), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n577), .A2(new_n584), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n572), .ZN(new_n975));
  OAI21_X1  g550(.A(G1981), .B1(new_n583), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n976), .A3(KEYINPUT49), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT49), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(new_n967), .A3(G8), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n967), .A2(G8), .A3(new_n968), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(KEYINPUT113), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n967), .A2(new_n985), .A3(G8), .A4(new_n968), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n949), .A2(new_n966), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2084), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n958), .A2(new_n989), .A3(new_n962), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n956), .B2(new_n957), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n924), .B1(new_n927), .B2(new_n926), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n753), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n958), .A2(new_n995), .A3(new_n962), .A4(new_n989), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(G8), .A3(G168), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n920), .B1(new_n988), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n964), .A2(new_n965), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n920), .ZN(new_n1001));
  INV_X1    g576(.A(new_n998), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n966), .A4(new_n987), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n983), .A2(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .A3(new_n986), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n972), .A2(new_n980), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n965), .A3(new_n964), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n934), .A2(new_n935), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n950), .B1(new_n1008), .B2(new_n924), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n980), .A2(new_n969), .A3(new_n779), .ZN(new_n1010));
  INV_X1    g585(.A(new_n974), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT115), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1007), .A2(new_n1015), .A3(new_n1012), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n999), .A2(new_n1003), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n991), .A2(G168), .A3(new_n994), .A4(new_n996), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n950), .A2(KEYINPUT124), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n997), .A2(G8), .A3(G286), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT62), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT51), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT62), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n1022), .A4(new_n1021), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n931), .A2(new_n932), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n697), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n958), .A2(new_n962), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1031), .A2(new_n1032), .B1(new_n798), .B2(new_n1033), .ZN(new_n1034));
  OR4_X1    g609(.A1(new_n1032), .A2(new_n992), .A3(G2078), .A4(new_n993), .ZN(new_n1035));
  AOI21_X1  g610(.A(G301), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n988), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1025), .A2(new_n1029), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(G1341), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n922), .A2(new_n924), .A3(new_n928), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT120), .B(G1996), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n967), .A2(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n548), .B1(new_n1044), .B2(KEYINPUT122), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n967), .A2(new_n1041), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1046), .A2(new_n1047), .A3(KEYINPUT122), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1039), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1348), .B1(new_n958), .B2(new_n962), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n967), .A2(G2067), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT60), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n598), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1956), .B1(new_n936), .B2(new_n943), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1042), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n558), .A2(new_n564), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  OR4_X1    g638(.A1(KEYINPUT61), .A2(new_n1057), .A3(new_n1059), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n939), .B1(new_n956), .B2(new_n957), .ZN(new_n1065));
  INV_X1    g640(.A(new_n942), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n924), .B1(new_n1066), .B2(new_n940), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n744), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1062), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1042), .A2(new_n1058), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(KEYINPUT61), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n1049), .A2(new_n1056), .A3(new_n1064), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1053), .A2(new_n598), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT118), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1068), .A2(new_n1081), .A3(new_n1071), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1063), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1080), .A2(new_n1082), .A3(KEYINPUT119), .A4(new_n1063), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n598), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1075), .A2(new_n1079), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n954), .A2(new_n829), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n821), .A2(new_n823), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1384), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT45), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(new_n1032), .A3(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n924), .A3(new_n922), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1033), .A2(new_n798), .ZN(new_n1097));
  AOI21_X1  g672(.A(G2078), .B1(new_n931), .B2(new_n932), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1096), .B(new_n1097), .C1(new_n1098), .C2(KEYINPUT53), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1090), .B1(new_n1036), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1027), .A2(new_n1022), .A3(new_n1021), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1034), .A2(G301), .A3(new_n1035), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(G171), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(KEYINPUT54), .A3(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1101), .A2(new_n1102), .A3(new_n1037), .A4(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1017), .B(new_n1038), .C1(new_n1089), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1094), .A2(new_n924), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT109), .ZN(new_n1109));
  INV_X1    g684(.A(G2067), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n716), .B(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1996), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1111), .B1(new_n726), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n938), .A2(new_n1093), .A3(KEYINPUT45), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(new_n1112), .A3(new_n726), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n769), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n767), .B(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(new_n1109), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G290), .B(G1986), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1107), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1115), .A2(new_n1112), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT46), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1109), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1111), .A2(new_n726), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT47), .Z(new_n1130));
  OR3_X1    g705(.A1(new_n1117), .A2(new_n1118), .A3(new_n767), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n717), .A2(new_n1110), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1108), .A2(G1986), .A3(G290), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT48), .Z(new_n1135));
  AOI211_X1 g710(.A(new_n1130), .B(new_n1133), .C1(new_n1120), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1124), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT125), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1124), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g716(.A1(G227), .A2(new_n465), .ZN(new_n1143));
  XOR2_X1   g717(.A(new_n1143), .B(KEYINPUT126), .Z(new_n1144));
  AND3_X1   g718(.A1(new_n1144), .A2(KEYINPUT127), .A3(new_n643), .ZN(new_n1145));
  AOI21_X1  g719(.A(KEYINPUT127), .B1(new_n1144), .B2(new_n643), .ZN(new_n1146));
  NOR3_X1   g720(.A1(G229), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g721(.A1(new_n916), .A2(new_n851), .A3(new_n1147), .ZN(G225));
  INV_X1    g722(.A(G225), .ZN(G308));
endmodule


