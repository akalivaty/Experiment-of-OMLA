//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  XOR2_X1   g002(.A(G127gat), .B(G134gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G141gat), .B(G148gat), .Z(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n211), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n205), .B(new_n215), .Z(new_n216));
  NAND2_X1  g015(.A1(G225gat), .A2(G233gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n205), .B1(KEYINPUT3), .B2(new_n215), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n213), .A2(new_n221), .A3(new_n214), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n217), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n225));
  INV_X1    g024(.A(new_n205), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(new_n215), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n215), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT77), .A3(new_n214), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n205), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n219), .B(KEYINPUT5), .C1(new_n224), .C2(new_n232), .ZN(new_n233));
  AOI211_X1 g032(.A(KEYINPUT5), .B(new_n218), .C1(new_n220), .C2(new_n222), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n226), .B2(new_n215), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(new_n225), .A3(new_n205), .A4(new_n230), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n234), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n234), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n233), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT0), .ZN(new_n243));
  XNOR2_X1  g042(.A(G57gat), .B(G85gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT6), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n233), .B(new_n248), .C1(new_n239), .C2(new_n240), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n245), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  NAND2_X1  g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n257), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G169gat), .ZN(new_n262));
  INV_X1    g061(.A(G176gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(KEYINPUT26), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n255), .A2(KEYINPUT71), .A3(new_n258), .A4(new_n256), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT27), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G183gat), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT27), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT69), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT28), .B(G190gat), .C1(new_n269), .C2(KEYINPUT68), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n279), .A2(new_n281), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G190gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(new_n284), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  AND2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n264), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(G169gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n287), .B1(new_n288), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n291), .A2(new_n296), .A3(KEYINPUT66), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT25), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n290), .A2(G169gat), .A3(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT67), .B1(new_n301), .B2(new_n289), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n256), .C1(new_n264), .C2(new_n290), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n264), .A2(new_n290), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT25), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n305), .A2(new_n287), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n283), .B1(new_n300), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(KEYINPUT75), .B(new_n283), .C1(new_n300), .C2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n313), .A2(new_n315), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319));
  INV_X1    g118(.A(G211gat), .ZN(new_n320));
  INV_X1    g119(.A(G218gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G211gat), .B(G218gat), .Z(new_n324));
  OR2_X1    g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n317), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n297), .A2(new_n288), .ZN(new_n330));
  INV_X1    g129(.A(new_n287), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n299), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n314), .B1(new_n336), .B2(new_n283), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n311), .A2(new_n338), .A3(new_n312), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n314), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(KEYINPUT76), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n342), .A3(new_n314), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n329), .B1(new_n344), .B2(new_n328), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n327), .B1(new_n341), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n329), .ZN(new_n353));
  INV_X1    g152(.A(new_n329), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n339), .A2(new_n342), .A3(new_n314), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n342), .B1(new_n339), .B2(new_n314), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n355), .A2(new_n356), .A3(new_n337), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n349), .C1(new_n357), .C2(new_n327), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n358), .A3(KEYINPUT30), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n253), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT64), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n205), .B1(new_n336), .B2(new_n283), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n205), .B(new_n283), .C1(new_n300), .C2(new_n308), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT33), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n366), .B2(KEYINPUT32), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n308), .B1(new_n333), .B2(new_n332), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n267), .A2(new_n278), .A3(new_n282), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n226), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n364), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT33), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n373), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n362), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n377), .B2(new_n364), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n370), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n385), .A2(KEYINPUT72), .A3(new_n379), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n372), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n382), .A3(new_n364), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n388), .B(KEYINPUT34), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n380), .A3(new_n373), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT72), .B1(new_n385), .B2(new_n379), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n389), .A3(new_n372), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n395), .A2(KEYINPUT74), .A3(new_n389), .A4(new_n372), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401));
  XNOR2_X1  g200(.A(G78gat), .B(G106gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT31), .B(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n327), .B1(new_n222), .B2(new_n338), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n230), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT77), .B1(new_n213), .B2(new_n214), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n325), .B2(new_n326), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n215), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT80), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n418), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n405), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n417), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(G22gat), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n416), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n405), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n401), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n416), .A2(new_n427), .ZN(new_n431));
  INV_X1    g230(.A(new_n426), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n404), .B1(new_n433), .B2(new_n423), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n434), .A2(new_n421), .A3(KEYINPUT81), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n360), .A2(new_n399), .A3(new_n400), .A4(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n436), .A2(new_n391), .A3(new_n396), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n438), .A2(new_n360), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(new_n400), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n238), .A2(new_n223), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n218), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(KEYINPUT39), .C1(new_n218), .C2(new_n216), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT39), .B(new_n217), .C1(new_n238), .C2(new_n223), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n444), .A2(new_n445), .A3(new_n245), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n447), .A3(new_n218), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT83), .B1(new_n448), .B2(new_n248), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT40), .B(new_n443), .C1(new_n446), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n246), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n444), .B2(new_n245), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n248), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT40), .B1(new_n454), .B2(new_n443), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n359), .A2(new_n456), .A3(new_n350), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(new_n436), .ZN(new_n458));
  NOR4_X1   g257(.A1(new_n355), .A2(new_n356), .A3(new_n328), .A4(new_n337), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n313), .A2(new_n315), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n309), .A2(new_n316), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n328), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n317), .A2(new_n464), .A3(new_n328), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n349), .B1(new_n345), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT85), .B(KEYINPUT37), .C1(new_n459), .C2(new_n466), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n354), .B1(new_n357), .B2(new_n327), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n351), .B1(new_n475), .B2(KEYINPUT37), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n345), .A2(new_n470), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n252), .B1(new_n345), .B2(new_n349), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n458), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n359), .A2(new_n350), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n252), .ZN(new_n483));
  INV_X1    g282(.A(new_n436), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n397), .A2(new_n398), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n391), .A2(KEYINPUT36), .A3(new_n396), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n483), .A2(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n481), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n483), .A2(new_n484), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n440), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(G197gat), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT11), .B(G169gat), .Z(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT12), .ZN(new_n500));
  AND2_X1   g299(.A1(G43gat), .A2(G50gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT15), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  INV_X1    g303(.A(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n506), .A2(KEYINPUT88), .A3(new_n507), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(KEYINPUT87), .C1(G29gat), .C2(G36gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT14), .ZN(new_n518));
  NOR3_X1   g317(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n514), .B(new_n516), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n516), .A2(new_n514), .ZN(new_n523));
  OR3_X1    g322(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(KEYINPUT14), .A3(new_n517), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n503), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n520), .B1(new_n512), .B2(new_n511), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT89), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n417), .A2(G15gat), .ZN(new_n533));
  INV_X1    g332(.A(G15gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n533), .B2(new_n535), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G1gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT92), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT91), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  OR3_X1    g342(.A1(new_n542), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n543), .B(new_n544), .C1(new_n537), .C2(new_n538), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n532), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547));
  INV_X1    g346(.A(new_n538), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  AND4_X1   g349(.A1(new_n547), .A2(new_n545), .A3(new_n550), .A4(new_n532), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n529), .B(new_n531), .C1(new_n546), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n529), .A2(new_n531), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n545), .A2(new_n550), .A3(new_n547), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G8gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n527), .A3(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n532), .A3(new_n545), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n552), .B(new_n553), .C1(new_n555), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT93), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n529), .A2(new_n531), .A3(new_n554), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n529), .A2(new_n531), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n559), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n564), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT18), .A4(new_n553), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n529), .A2(new_n531), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n557), .A3(new_n559), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n552), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n553), .B(KEYINPUT13), .Z(new_n575));
  AOI22_X1  g374(.A1(new_n561), .A2(new_n562), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n500), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n500), .ZN(new_n580));
  AOI211_X1 g379(.A(KEYINPUT86), .B(new_n580), .C1(new_n571), .C2(new_n576), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT10), .ZN(new_n584));
  INV_X1    g383(.A(G57gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT94), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G57gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n588), .A3(G64gat), .ZN(new_n589));
  INV_X1    g388(.A(G64gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G57gat), .ZN(new_n591));
  AND2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT9), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n589), .A2(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n585), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(KEYINPUT9), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT95), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n592), .A2(new_n594), .ZN(new_n603));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n591), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(G57gat), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(G64gat), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n592), .B1(KEYINPUT9), .B2(new_n594), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n602), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(KEYINPUT98), .A2(G99gat), .A3(G106gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT8), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g415(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT99), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n616), .A2(new_n619), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n616), .A2(new_n619), .A3(new_n625), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n601), .A2(new_n611), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n632), .A2(new_n630), .A3(new_n627), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n584), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n627), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n601), .A2(new_n611), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT10), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OR3_X1    g440(.A1(new_n631), .A2(new_n633), .A3(new_n640), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  OR2_X1    g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n583), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n567), .B1(KEYINPUT21), .B2(new_n637), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT96), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n655), .B(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n565), .A2(new_n558), .A3(new_n635), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n566), .A2(new_n636), .ZN(new_n665));
  XNOR2_X1  g464(.A(G190gat), .B(G218gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  AND2_X1   g466(.A1(G232gat), .A2(G233gat), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n667), .A2(KEYINPUT101), .B1(KEYINPUT41), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G134gat), .B(G162gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n668), .A2(KEYINPUT41), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n671), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n664), .A2(new_n665), .A3(new_n669), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n672), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n672), .B2(new_n677), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n650), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n252), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n540), .ZN(G1324gat));
  INV_X1    g485(.A(new_n684), .ZN(new_n687));
  INV_X1    g486(.A(new_n482), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n532), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n684), .A2(new_n482), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n493), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n487), .A2(KEYINPUT102), .A3(new_n488), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n684), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n399), .A2(new_n534), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n684), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n436), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n650), .A2(new_n663), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n495), .A2(new_n681), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(G29gat), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n707), .A3(new_n253), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n481), .A2(new_n695), .A3(new_n492), .A4(new_n696), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n440), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n679), .B2(new_n680), .ZN(new_n713));
  INV_X1    g512(.A(new_n680), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT103), .A3(new_n678), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n681), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n492), .A2(new_n493), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT82), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n489), .A2(new_n490), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n481), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(new_n440), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n705), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n253), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n709), .B1(new_n728), .B2(new_n707), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n706), .A2(new_n730), .A3(new_n688), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n726), .A2(new_n688), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(new_n730), .ZN(G1329gat));
  INV_X1    g535(.A(new_n697), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n724), .B1(new_n495), .B2(new_n681), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n711), .A2(new_n716), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n737), .B(new_n705), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n706), .A2(new_n504), .A3(new_n399), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1330gat));
  NAND4_X1  g545(.A1(new_n495), .A2(KEYINPUT104), .A3(new_n681), .A4(new_n705), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n484), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT104), .B1(new_n723), .B2(new_n705), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n505), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n725), .A2(G50gat), .A3(new_n484), .A4(new_n705), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n750), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1331gat));
  NAND3_X1  g555(.A1(new_n583), .A2(new_n649), .A3(new_n682), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n710), .B2(new_n440), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n253), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(new_n608), .Z(G1332gat));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n688), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT49), .B(G64gat), .Z(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(G1333gat));
  XOR2_X1   g563(.A(new_n399), .B(KEYINPUT105), .Z(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(G71gat), .B1(new_n758), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n737), .A2(G71gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n484), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n621), .A2(new_n623), .ZN(new_n773));
  INV_X1    g572(.A(new_n649), .ZN(new_n774));
  INV_X1    g573(.A(new_n663), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n582), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n725), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n777), .B2(new_n252), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n582), .A2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n681), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n711), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n783), .B(new_n780), .C1(new_n710), .C2(new_n440), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n252), .A2(new_n773), .A3(new_n774), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT106), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n786), .B2(new_n788), .ZN(G1336gat));
  OAI211_X1 g588(.A(new_n688), .B(new_n776), .C1(new_n738), .C2(new_n739), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT107), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n725), .A2(new_n792), .A3(new_n688), .A4(new_n776), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(G92gat), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n482), .A2(G92gat), .A3(new_n774), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n790), .A2(G92gat), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n785), .A2(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n777), .B2(new_n697), .ZN(new_n802));
  INV_X1    g601(.A(G99gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n399), .A2(new_n803), .A3(new_n649), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n786), .B2(new_n804), .ZN(G1338gat));
  OAI211_X1 g604(.A(new_n484), .B(new_n776), .C1(new_n738), .C2(new_n739), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n725), .A2(KEYINPUT109), .A3(new_n484), .A4(new_n776), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(G106gat), .A3(new_n809), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n436), .A2(G106gat), .A3(new_n774), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n782), .B2(new_n784), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT108), .B(new_n811), .C1(new_n782), .C2(new_n784), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n806), .A2(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n812), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n713), .A2(new_n715), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n639), .B2(new_n640), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n827));
  INV_X1    g626(.A(new_n640), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n634), .A2(new_n827), .A3(new_n828), .A4(new_n638), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n634), .A2(new_n828), .A3(new_n638), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT110), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n634), .B2(new_n638), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n646), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n824), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n832), .C2(new_n834), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n836), .B(new_n646), .C1(new_n833), .C2(new_n825), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n832), .A3(KEYINPUT111), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n648), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT111), .B1(new_n840), .B2(new_n832), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n561), .A2(new_n562), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n574), .A2(new_n575), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n563), .B2(new_n570), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n580), .B1(new_n848), .B2(KEYINPUT86), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n577), .A2(new_n578), .A3(new_n500), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n839), .A2(new_n844), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n571), .A2(new_n576), .A3(new_n500), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n568), .A2(new_n553), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n574), .A2(new_n575), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n499), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n649), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n823), .B1(new_n851), .B2(new_n858), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n823), .A2(new_n857), .A3(new_n844), .A4(new_n839), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n822), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n826), .A2(new_n829), .A3(new_n831), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n834), .A2(KEYINPUT55), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n648), .A3(new_n841), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n837), .A3(new_n838), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n823), .A3(new_n857), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n774), .A2(new_n856), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n867), .B2(new_n582), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT113), .B(new_n868), .C1(new_n870), .C2(new_n823), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n861), .A2(new_n871), .A3(new_n663), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n583), .A2(new_n774), .A3(new_n682), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n484), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n688), .A2(new_n252), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n399), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(G113gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n583), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n252), .B1(new_n872), .B2(new_n873), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n438), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n482), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n582), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n885), .B2(new_n878), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n887), .A3(new_n649), .ZN(new_n888));
  OAI21_X1  g687(.A(G120gat), .B1(new_n877), .B2(new_n774), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n893), .A3(new_n775), .ZN(new_n894));
  OAI21_X1  g693(.A(G127gat), .B1(new_n877), .B2(new_n663), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1342gat));
  NOR2_X1   g695(.A1(new_n718), .A2(G134gat), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n482), .A3(new_n883), .A4(new_n897), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n877), .B2(new_n718), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT116), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n898), .B2(KEYINPUT56), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n899), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(G1343gat));
  NOR3_X1   g704(.A1(new_n737), .A2(new_n688), .A3(new_n436), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n583), .A2(G141gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n880), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT58), .B1(new_n908), .B2(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n697), .A2(new_n875), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n872), .A2(new_n873), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n484), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n484), .A2(KEYINPUT57), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n835), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n582), .A2(new_n844), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n681), .B1(new_n917), .B2(new_n858), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n663), .B1(new_n918), .B2(new_n860), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n914), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n911), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G141gat), .B1(new_n921), .B2(new_n583), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n909), .B(new_n922), .C1(KEYINPUT120), .C2(new_n908), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n925), .B(new_n911), .C1(new_n913), .C2(new_n920), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n582), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n906), .A2(new_n880), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n927), .A2(G141gat), .B1(new_n928), .B2(new_n907), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(G1344gat));
  NAND3_X1  g730(.A1(new_n912), .A2(KEYINPUT57), .A3(new_n484), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n867), .A2(new_n681), .A3(new_n857), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n663), .B1(new_n918), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n436), .B1(new_n934), .B2(new_n873), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(KEYINPUT57), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n774), .B1(new_n910), .B2(KEYINPUT121), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(new_n937), .C1(KEYINPUT121), .C2(new_n910), .ZN(new_n938));
  AND2_X1   g737(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n774), .A2(G148gat), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(new_n928), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n649), .A3(new_n926), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(G148gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n943), .B2(KEYINPUT59), .ZN(G1345gat));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n926), .ZN(new_n945));
  OAI21_X1  g744(.A(G155gat), .B1(new_n945), .B2(new_n663), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n207), .A3(new_n775), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1346gat));
  NAND3_X1  g747(.A1(new_n924), .A2(new_n823), .A3(new_n926), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n924), .A2(KEYINPUT122), .A3(new_n823), .A4(new_n926), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(G162gat), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n928), .A2(new_n208), .A3(new_n681), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n482), .A2(new_n253), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n874), .A2(new_n766), .A3(new_n956), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(new_n262), .A3(new_n583), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n912), .A2(new_n438), .A3(new_n956), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n582), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n958), .A2(new_n960), .ZN(G1348gat));
  AOI21_X1  g760(.A(G176gat), .B1(new_n959), .B2(new_n649), .ZN(new_n962));
  INV_X1    g761(.A(new_n957), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n774), .B1(new_n293), .B2(new_n295), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1349gat));
  AND3_X1   g764(.A1(new_n775), .A2(new_n273), .A3(new_n276), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n963), .A2(new_n775), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(G183gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT60), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n968), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n274), .A3(new_n823), .ZN(new_n977));
  OAI21_X1  g776(.A(G190gat), .B1(new_n957), .B2(new_n718), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(G1351gat));
  AND2_X1   g783(.A1(new_n697), .A2(new_n956), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n985), .A2(new_n484), .A3(new_n912), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n582), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n936), .A2(new_n985), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n582), .A2(G197gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  XNOR2_X1  g791(.A(KEYINPUT126), .B(G204gat), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n986), .A2(new_n774), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n993), .B1(new_n989), .B2(new_n774), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1353gat));
  NAND3_X1  g796(.A1(new_n987), .A2(new_n320), .A3(new_n775), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n936), .A2(new_n775), .A3(new_n985), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n999), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT63), .B1(new_n999), .B2(G211gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n989), .B2(new_n718), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n321), .A3(new_n823), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1003), .A2(KEYINPUT127), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


