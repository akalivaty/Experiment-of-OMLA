//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946;
  XNOR2_X1  g000(.A(G169gat), .B(G197gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT85), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G113gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT86), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n203), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n206), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT12), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n208), .A2(new_n213), .A3(KEYINPUT12), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT13), .ZN(new_n220));
  INV_X1    g019(.A(G22gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G15gat), .ZN(new_n222));
  INV_X1    g021(.A(G15gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G22gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(KEYINPUT88), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(KEYINPUT88), .B2(new_n226), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n231));
  XNOR2_X1  g030(.A(G15gat), .B(G22gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G8gat), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT89), .B1(new_n225), .B2(new_n226), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n229), .A2(new_n227), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n235), .B(new_n236), .C1(new_n237), .C2(new_n225), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G29gat), .A2(G36gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G50gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G43gat), .ZN(new_n246));
  INV_X1    g045(.A(G43gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G50gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT15), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(G50gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n245), .A2(G43gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(new_n240), .A3(new_n249), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n257));
  INV_X1    g056(.A(G29gat), .ZN(new_n258));
  INV_X1    g057(.A(G36gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT87), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n259), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n242), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n251), .B1(new_n256), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n239), .A2(new_n266), .ZN(new_n267));
  NOR4_X1   g066(.A1(KEYINPUT87), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n263), .B1(new_n262), .B2(new_n259), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n241), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G43gat), .B(G50gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n255), .A3(new_n272), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n234), .A2(new_n238), .B1(new_n273), .B2(new_n251), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n220), .B1(new_n267), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n234), .A2(new_n238), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT17), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n251), .B(new_n278), .C1(new_n256), .C2(new_n265), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n273), .B2(new_n251), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n219), .A3(new_n275), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT18), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n266), .A2(KEYINPUT17), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n239), .B1(new_n287), .B2(new_n279), .ZN(new_n288));
  INV_X1    g087(.A(new_n219), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n288), .A2(new_n289), .A3(new_n274), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n286), .B1(new_n290), .B2(KEYINPUT18), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n282), .A2(KEYINPUT18), .A3(new_n219), .A4(new_n275), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT90), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n218), .B(new_n285), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT91), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n292), .B(KEYINPUT90), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n297), .A2(KEYINPUT91), .A3(new_n218), .A4(new_n285), .ZN(new_n298));
  INV_X1    g097(.A(new_n218), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n285), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n296), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT23), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n304), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n318), .A2(new_n304), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n308), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(new_n306), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n319), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n308), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n312), .A2(KEYINPUT26), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n317), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT65), .A2(KEYINPUT26), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT65), .A2(KEYINPUT26), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n315), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(KEYINPUT66), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n325), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT1), .ZN(new_n342));
  XOR2_X1   g141(.A(G127gat), .B(G134gat), .Z(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n303), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n339), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n308), .A3(new_n330), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n348), .A2(KEYINPUT67), .A3(new_n344), .A4(new_n325), .ZN(new_n349));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n340), .A2(new_n345), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n346), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT34), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(KEYINPUT34), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n356));
  INV_X1    g155(.A(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G15gat), .B(G43gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G71gat), .B(G99gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(new_n356), .B2(new_n357), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT33), .B1(new_n356), .B2(new_n357), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n302), .B(new_n355), .C1(new_n365), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n355), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n370), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(KEYINPUT68), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT36), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT69), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n353), .A2(KEYINPUT69), .A3(new_n354), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT36), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n376), .A3(new_n355), .A4(new_n370), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(KEYINPUT70), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G141gat), .B(G148gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(G155gat), .B2(G162gat), .ZN(new_n386));
  AND2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387));
  OAI22_X1  g186(.A1(new_n384), .A2(new_n386), .B1(KEYINPUT74), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G155gat), .B(G162gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n388), .B(new_n389), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n344), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n345), .B2(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n344), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n401));
  OR3_X1    g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT5), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n400), .B2(KEYINPUT5), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n345), .B(new_n393), .ZN(new_n405));
  INV_X1    g204(.A(new_n398), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n402), .A2(new_n403), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT6), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(KEYINPUT79), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n400), .ZN(new_n417));
  INV_X1    g216(.A(new_n403), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT5), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n408), .A2(KEYINPUT83), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT72), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n340), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n432), .B(KEYINPUT71), .Z(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n348), .B2(new_n325), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G197gat), .B(G204gat), .Z(new_n437));
  AOI21_X1  g236(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G211gat), .B(G218gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n434), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n441), .ZN(new_n443));
  INV_X1    g242(.A(new_n433), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n340), .B2(new_n430), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n445), .B2(new_n435), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n429), .B1(new_n447), .B2(KEYINPUT37), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT38), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n442), .A2(new_n429), .A3(new_n446), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n448), .A2(new_n451), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n413), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n424), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT80), .B(KEYINPUT39), .Z(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n406), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n415), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT81), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n465), .A3(new_n415), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n406), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(KEYINPUT39), .C1(new_n406), .C2(new_n405), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n415), .B1(new_n408), .B2(KEYINPUT83), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n420), .A2(new_n421), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n447), .A2(new_n428), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n442), .A2(new_n446), .A3(KEYINPUT30), .A4(new_n429), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n469), .A2(new_n470), .A3(new_n459), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n472), .A2(new_n475), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n484), .B(KEYINPUT78), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G78gat), .B(G106gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT31), .B(G50gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n221), .ZN(new_n490));
  NAND2_X1  g289(.A1(KEYINPUT77), .A2(G22gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n489), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n441), .B1(new_n392), .B2(new_n430), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n441), .A2(new_n430), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n390), .B1(new_n494), .B2(new_n391), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n493), .A2(new_n495), .A3(new_n492), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n486), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n485), .A3(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n458), .A2(new_n483), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n420), .B2(new_n456), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n408), .A2(new_n413), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n457), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n476), .A2(new_n477), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT73), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n476), .A2(KEYINPUT73), .A3(new_n477), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(new_n480), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n502), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n383), .A2(new_n503), .A3(new_n504), .A4(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n502), .B1(new_n371), .B2(new_n374), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT35), .B1(new_n518), .B2(new_n514), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n478), .A2(new_n520), .A3(new_n502), .A4(new_n480), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n379), .B2(new_n381), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n424), .A2(new_n457), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n301), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G78gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G64gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G57gat), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n535));
  INV_X1    g334(.A(G57gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G64gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT92), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT93), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n532), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n277), .B1(new_n527), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n527), .ZN(new_n545));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT94), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n548), .B(new_n554), .Z(new_n555));
  XNOR2_X1  g354(.A(G99gat), .B(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT96), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(G85gat), .A3(G92gat), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n557), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT7), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n556), .A3(new_n564), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(KEYINPUT97), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n562), .A2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n556), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n266), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n280), .A2(new_n281), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n583), .A2(new_n584), .B1(new_n585), .B2(new_n579), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT99), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n586), .A2(new_n588), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n589), .A2(new_n595), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n592), .B(KEYINPUT100), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n575), .A2(new_n578), .A3(new_n542), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n540), .B(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(new_n528), .A3(new_n538), .A4(new_n535), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n532), .A3(new_n574), .A4(new_n571), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n601), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT101), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n602), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n532), .B(KEYINPUT10), .C1(new_n539), .C2(new_n541), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n579), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n601), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n608), .A2(new_n619), .A3(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n555), .A2(new_n600), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n526), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n508), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT102), .B(G1gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1324gat));
  INV_X1    g429(.A(new_n481), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n228), .A2(new_n236), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n236), .B2(new_n632), .ZN(new_n636));
  MUX2_X1   g435(.A(new_n635), .B(new_n636), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g436(.A1(new_n379), .A2(new_n381), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n223), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n383), .A2(new_n504), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(new_n627), .A3(new_n223), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n641), .A2(new_n647), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n526), .A2(new_n515), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n625), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT105), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT43), .B(G22gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  AOI21_X1  g452(.A(new_n600), .B1(new_n517), .B2(new_n525), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n555), .A2(new_n301), .A3(new_n623), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n508), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n258), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT106), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT45), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n661));
  AOI221_X4 g460(.A(new_n366), .B1(KEYINPUT33), .B2(new_n364), .C1(new_n356), .C2(new_n357), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT68), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n355), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n373), .A2(KEYINPUT68), .A3(new_n372), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n515), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n511), .A2(new_n512), .A3(new_n480), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n420), .A2(new_n456), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n414), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n669), .B2(new_n457), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n520), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n522), .A2(new_n523), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT107), .B1(new_n519), .B2(new_n524), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n517), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n599), .B1(new_n589), .B2(new_n595), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n594), .B2(new_n597), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n676), .A2(new_n677), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n673), .B1(new_n671), .B2(new_n672), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n519), .A2(KEYINPUT107), .A3(new_n524), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n382), .A2(KEYINPUT70), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n375), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n469), .A2(new_n470), .A3(new_n459), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n471), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n473), .A2(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n515), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n690), .A2(new_n458), .B1(new_n515), .B2(new_n514), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n682), .A2(new_n683), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n600), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT108), .B1(new_n654), .B2(new_n678), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n655), .B(new_n681), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n508), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n660), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n656), .A2(new_n259), .A3(new_n481), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  NOR2_X1   g498(.A1(new_n695), .A2(new_n631), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n700), .B2(KEYINPUT109), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  OAI21_X1  g503(.A(G43gat), .B1(new_n695), .B2(new_n686), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n639), .A2(G43gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n656), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n704), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n517), .A2(new_n525), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n680), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n713), .A3(KEYINPUT108), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n714), .A2(new_n645), .A3(new_n655), .A4(new_n681), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n709), .B1(new_n715), .B2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT110), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G43gat), .B1(new_n695), .B2(new_n646), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n704), .A3(new_n707), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n714), .A2(new_n642), .A3(new_n655), .A4(new_n681), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(G43gat), .B1(new_n656), .B2(new_n706), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n719), .B(new_n720), .C1(new_n704), .C2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n717), .A2(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n695), .B2(new_n502), .ZN(new_n725));
  INV_X1    g524(.A(new_n555), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n726), .A2(new_n245), .A3(new_n680), .A4(new_n624), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n649), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g528(.A1(new_n296), .A2(new_n298), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n300), .A2(new_n299), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n555), .A2(new_n600), .A3(new_n623), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n692), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n657), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n481), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n734), .A2(new_n645), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n639), .A2(G71gat), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(G71gat), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n515), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT111), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  NOR2_X1   g546(.A1(new_n555), .A2(new_n732), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n714), .A2(new_n623), .A3(new_n681), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n508), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n692), .A2(new_n600), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n748), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n751), .A2(new_n748), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n754), .A2(KEYINPUT113), .A3(new_n755), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n623), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n657), .A2(new_n567), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n750), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n749), .B2(new_n631), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n631), .A2(G92gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n623), .B(new_n764), .C1(new_n754), .C2(new_n755), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT52), .ZN(G1337gat));
  XNOR2_X1  g566(.A(KEYINPUT114), .B(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n749), .B2(new_n646), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n639), .A2(new_n768), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n760), .B2(new_n770), .ZN(G1338gat));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n502), .A2(G106gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n623), .B(new_n773), .C1(new_n754), .C2(new_n755), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(KEYINPUT115), .ZN(new_n775));
  OAI21_X1  g574(.A(G106gat), .B1(new_n749), .B2(new_n502), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n774), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n775), .B(new_n777), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  INV_X1    g579(.A(new_n601), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n610), .B2(new_n613), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n780), .B(new_n619), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n601), .B1(new_n579), .B2(new_n612), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n610), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT54), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(KEYINPUT116), .A3(new_n782), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n783), .B1(new_n610), .B2(new_n785), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n615), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n784), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n622), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT116), .B1(new_n787), .B2(new_n782), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n615), .A2(new_n789), .A3(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n619), .B1(new_n782), .B2(new_n783), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n732), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n289), .B1(new_n288), .B2(new_n274), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n267), .A2(new_n275), .A3(new_n220), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n214), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n296), .B2(new_n298), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n623), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n680), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n680), .A2(new_n804), .A3(new_n799), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n779), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n680), .A2(new_n799), .A3(new_n804), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n732), .A2(new_n799), .B1(new_n804), .B2(new_n623), .ZN(new_n810));
  OAI211_X1 g609(.A(KEYINPUT117), .B(new_n809), .C1(new_n810), .C2(new_n680), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n726), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n625), .A2(new_n732), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n817), .A3(new_n515), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n657), .A3(new_n638), .A4(new_n631), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n209), .A3(new_n301), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n816), .A2(new_n817), .A3(new_n508), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n518), .A2(new_n481), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n732), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n209), .B2(new_n823), .ZN(G1340gat));
  INV_X1    g623(.A(G120gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n819), .A2(new_n825), .A3(new_n624), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n623), .A3(new_n822), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(G1341gat));
  OAI21_X1  g627(.A(G127gat), .B1(new_n819), .B2(new_n726), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n821), .A2(new_n822), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n726), .A2(G127gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G1342gat));
  OR2_X1    g631(.A1(new_n819), .A2(new_n600), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n830), .A2(G134gat), .A3(new_n600), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n833), .A2(G134gat), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(G1343gat));
  NAND3_X1  g640(.A1(new_n686), .A2(new_n657), .A3(new_n631), .ZN(new_n842));
  INV_X1    g641(.A(new_n805), .ZN(new_n843));
  INV_X1    g642(.A(new_n797), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n794), .B2(new_n795), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n622), .B(new_n792), .C1(new_n845), .C2(KEYINPUT55), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n301), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n600), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n807), .B1(new_n848), .B2(KEYINPUT120), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n555), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n515), .B1(new_n851), .B2(new_n814), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n842), .B1(new_n852), .B2(KEYINPUT57), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n812), .A2(new_n815), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n515), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n211), .B1(new_n859), .B2(new_n732), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n481), .A2(new_n502), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n646), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(G141gat), .A3(new_n301), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n860), .B2(KEYINPUT121), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n864), .B(new_n866), .ZN(G1344gat));
  OR3_X1    g666(.A1(new_n862), .A2(G148gat), .A3(new_n624), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n855), .A2(new_n515), .A3(new_n857), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n555), .B1(new_n848), .B2(new_n809), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n856), .B(new_n515), .C1(new_n872), .C2(new_n814), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n842), .A2(new_n624), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n869), .A2(G148gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n859), .B2(new_n623), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n868), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1345gat));
  INV_X1    g680(.A(new_n859), .ZN(new_n882));
  OAI21_X1  g681(.A(G155gat), .B1(new_n882), .B2(new_n726), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n726), .A2(G155gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n862), .B2(new_n884), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n859), .A2(G162gat), .A3(new_n680), .ZN(new_n886));
  INV_X1    g685(.A(G162gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n862), .B2(new_n600), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n657), .A2(new_n631), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR4_X1   g690(.A1(new_n816), .A2(new_n817), .A3(new_n518), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n310), .A3(new_n732), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT123), .Z(new_n894));
  NAND3_X1  g693(.A1(new_n818), .A2(new_n638), .A3(new_n890), .ZN(new_n895));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n301), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1348gat));
  OAI21_X1  g696(.A(G176gat), .B1(new_n895), .B2(new_n624), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n311), .A3(new_n623), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1349gat));
  OAI21_X1  g699(.A(G183gat), .B1(new_n895), .B2(new_n726), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n892), .A2(new_n326), .A3(new_n555), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n892), .A2(new_n327), .A3(new_n680), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n895), .A2(new_n600), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  NOR2_X1   g710(.A1(new_n645), .A2(new_n891), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n816), .A2(new_n817), .A3(new_n502), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n873), .B(new_n912), .C1(new_n913), .C2(new_n856), .ZN(new_n914));
  INV_X1    g713(.A(G197gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n301), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n912), .A3(new_n732), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n913), .A2(new_n912), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n624), .A2(G204gat), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  OAI21_X1  g723(.A(G204gat), .B1(new_n914), .B2(new_n624), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G1353gat));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n914), .A2(new_n726), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n930));
  INV_X1    g729(.A(G211gat), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(KEYINPUT125), .B2(new_n932), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n929), .A2(new_n933), .B1(new_n928), .B2(KEYINPUT63), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n555), .A2(new_n931), .ZN(new_n935));
  OAI22_X1  g734(.A1(new_n930), .A2(new_n934), .B1(new_n919), .B2(new_n935), .ZN(G1354gat));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n914), .A2(KEYINPUT126), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n871), .A2(new_n939), .A3(new_n873), .A4(new_n912), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n680), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G218gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n919), .A2(G218gat), .A3(new_n600), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n937), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g744(.A(KEYINPUT127), .B(new_n943), .C1(new_n941), .C2(G218gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1355gat));
endmodule


