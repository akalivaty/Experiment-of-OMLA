

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XOR2_X1 U321 ( .A(G22GAT), .B(G155GAT), .Z(n431) );
  XNOR2_X1 U322 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U323 ( .A(n333), .B(n332), .ZN(n335) );
  XNOR2_X1 U324 ( .A(n388), .B(n387), .ZN(n526) );
  XNOR2_X1 U325 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n404) );
  XNOR2_X1 U326 ( .A(n405), .B(n404), .ZN(n563) );
  XOR2_X1 U327 ( .A(n342), .B(n372), .Z(n482) );
  NOR2_X1 U328 ( .A1(n527), .A2(n447), .ZN(n556) );
  XOR2_X1 U329 ( .A(n568), .B(KEYINPUT41), .Z(n545) );
  XOR2_X1 U330 ( .A(n464), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U331 ( .A(n448), .B(G190GAT), .ZN(n449) );
  XNOR2_X1 U332 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U333 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G127GAT), .B(G134GAT), .Z(n290) );
  XNOR2_X1 U335 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U337 ( .A(G113GAT), .B(n291), .Z(n427) );
  XOR2_X1 U338 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U339 ( .A(G71GAT), .B(G176GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n427), .B(n294), .ZN(n306) );
  XOR2_X1 U342 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n296) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n399) );
  XOR2_X1 U345 ( .A(G190GAT), .B(n399), .Z(n298) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U348 ( .A(G183GAT), .B(KEYINPUT84), .Z(n300) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U351 ( .A(n302), .B(n301), .Z(n304) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n527) );
  XOR2_X1 U355 ( .A(KEYINPUT66), .B(KEYINPUT76), .Z(n308) );
  XNOR2_X1 U356 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  XOR2_X1 U359 ( .A(n309), .B(n361), .Z(n311) );
  XNOR2_X1 U360 ( .A(G218GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U362 ( .A(n312), .B(KEYINPUT77), .Z(n316) );
  XOR2_X1 U363 ( .A(G29GAT), .B(G43GAT), .Z(n314) );
  XNOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n350) );
  XNOR2_X1 U366 ( .A(n350), .B(G134GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n325) );
  XOR2_X1 U368 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n318) );
  XNOR2_X1 U369 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U371 ( .A(G36GAT), .B(G190GAT), .Z(n394) );
  XNOR2_X1 U372 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n319), .B(G162GAT), .ZN(n435) );
  XOR2_X1 U374 ( .A(n394), .B(n435), .Z(n321) );
  NAND2_X1 U375 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U377 ( .A(n323), .B(n322), .Z(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n552) );
  XOR2_X1 U379 ( .A(KEYINPUT15), .B(n431), .Z(n327) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U381 ( .A(n353), .B(G127GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n329) );
  XNOR2_X1 U384 ( .A(KEYINPUT80), .B(KEYINPUT12), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n331) );
  AND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  INV_X1 U387 ( .A(KEYINPUT14), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n338) );
  XNOR2_X1 U389 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(G211GAT), .ZN(n397) );
  XNOR2_X1 U391 ( .A(G64GAT), .B(n397), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .Z(n340) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(G78GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT68), .B(n341), .Z(n372) );
  INV_X1 U397 ( .A(n482), .ZN(n343) );
  XOR2_X1 U398 ( .A(n343), .B(KEYINPUT111), .Z(n557) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G22GAT), .Z(n345) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G197GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n347) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(G8GAT), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n358) );
  XOR2_X1 U406 ( .A(n350), .B(KEYINPUT29), .Z(n352) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n356) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n564) );
  XOR2_X1 U413 ( .A(G64GAT), .B(G92GAT), .Z(n360) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(G204GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n400) );
  XOR2_X1 U416 ( .A(KEYINPUT32), .B(n400), .Z(n363) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n368) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n364), .B(G148GAT), .ZN(n438) );
  XOR2_X1 U421 ( .A(n438), .B(KEYINPUT31), .Z(n366) );
  NAND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n365) );
  XOR2_X1 U423 ( .A(n366), .B(n365), .Z(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n374) );
  XOR2_X1 U425 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n370) );
  XNOR2_X1 U426 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n568) );
  NAND2_X1 U430 ( .A1(n564), .A2(n545), .ZN(n375) );
  XOR2_X1 U431 ( .A(n375), .B(KEYINPUT46), .Z(n376) );
  NOR2_X1 U432 ( .A1(n557), .A2(n376), .ZN(n377) );
  XOR2_X1 U433 ( .A(KEYINPUT112), .B(n377), .Z(n378) );
  NOR2_X1 U434 ( .A1(n552), .A2(n378), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n379), .B(KEYINPUT47), .ZN(n386) );
  XOR2_X1 U436 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n382) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n380), .B(n552), .ZN(n576) );
  NOR2_X1 U439 ( .A1(n576), .A2(n482), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n383) );
  NOR2_X1 U441 ( .A1(n568), .A2(n383), .ZN(n384) );
  INV_X1 U442 ( .A(n564), .ZN(n497) );
  NAND2_X1 U443 ( .A1(n384), .A2(n497), .ZN(n385) );
  NAND2_X1 U444 ( .A1(n386), .A2(n385), .ZN(n388) );
  XNOR2_X1 U445 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n387) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n390) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(G218GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n440) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(n440), .Z(n392) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U452 ( .A(n393), .B(KEYINPUT94), .Z(n396) );
  XNOR2_X1 U453 ( .A(n394), .B(KEYINPUT93), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U455 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U457 ( .A(n402), .B(n401), .Z(n515) );
  INV_X1 U458 ( .A(n515), .ZN(n403) );
  NAND2_X1 U459 ( .A1(n526), .A2(n403), .ZN(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT89), .B(KEYINPUT92), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G155GAT), .Z(n409) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(G148GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U466 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(G141GAT), .B(n414), .Z(n441) );
  XOR2_X1 U471 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n416) );
  XNOR2_X1 U472 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n441), .B(n417), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U476 ( .A(KEYINPUT88), .B(KEYINPUT6), .Z(n421) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U479 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n561) );
  XOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n429) );
  XNOR2_X1 U484 ( .A(KEYINPUT23), .B(G78GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U486 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U489 ( .A(n434), .B(G204GAT), .Z(n437) );
  XNOR2_X1 U490 ( .A(n435), .B(G211GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n464) );
  INV_X1 U495 ( .A(n464), .ZN(n444) );
  AND2_X1 U496 ( .A1(n561), .A2(n444), .ZN(n445) );
  AND2_X1 U497 ( .A1(n563), .A2(n445), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n556), .A2(n552), .ZN(n450) );
  XOR2_X1 U500 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n448) );
  NAND2_X1 U501 ( .A1(n556), .A2(n545), .ZN(n456) );
  XOR2_X1 U502 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n452) );
  XNOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(n454) );
  XOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT122), .Z(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NOR2_X1 U508 ( .A1(n568), .A2(n497), .ZN(n457) );
  XOR2_X1 U509 ( .A(KEYINPUT73), .B(n457), .Z(n486) );
  XNOR2_X1 U510 ( .A(n515), .B(KEYINPUT27), .ZN(n524) );
  NAND2_X1 U511 ( .A1(n529), .A2(n527), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n524), .A2(n458), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n561), .A2(n459), .ZN(n469) );
  NOR2_X1 U514 ( .A1(n527), .A2(n515), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n464), .A2(n460), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT96), .B(n461), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT25), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n463), .A2(n561), .ZN(n467) );
  NAND2_X1 U519 ( .A1(n464), .A2(n527), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT26), .ZN(n559) );
  NOR2_X1 U521 ( .A1(n524), .A2(n559), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n484) );
  NOR2_X1 U524 ( .A1(n482), .A2(n552), .ZN(n470) );
  XOR2_X1 U525 ( .A(KEYINPUT81), .B(n470), .Z(n471) );
  XNOR2_X1 U526 ( .A(KEYINPUT16), .B(n471), .ZN(n472) );
  AND2_X1 U527 ( .A1(n484), .A2(n472), .ZN(n499) );
  NAND2_X1 U528 ( .A1(n486), .A2(n499), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n561), .A2(n479), .ZN(n473) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n473), .Z(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(n474), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n515), .A2(n479), .ZN(n475) );
  XOR2_X1 U533 ( .A(G8GAT), .B(n475), .Z(G1325GAT) );
  NOR2_X1 U534 ( .A1(n527), .A2(n479), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT35), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U537 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NOR2_X1 U538 ( .A1(n529), .A2(n479), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(n480), .Z(n481) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U541 ( .A1(n576), .A2(n343), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n485), .ZN(n512) );
  NAND2_X1 U544 ( .A1(n512), .A2(n486), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n495) );
  NOR2_X1 U547 ( .A1(n561), .A2(n495), .ZN(n490) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n515), .A2(n495), .ZN(n491) );
  XOR2_X1 U551 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U552 ( .A1(n527), .A2(n495), .ZN(n493) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U556 ( .A1(n529), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  NAND2_X1 U558 ( .A1(n497), .A2(n545), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(KEYINPUT103), .ZN(n511) );
  NAND2_X1 U560 ( .A1(n511), .A2(n499), .ZN(n505) );
  NOR2_X1 U561 ( .A1(n561), .A2(n505), .ZN(n501) );
  XNOR2_X1 U562 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U565 ( .A1(n515), .A2(n505), .ZN(n503) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n527), .A2(n505), .ZN(n504) );
  XOR2_X1 U568 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U569 ( .A1(n529), .A2(n505), .ZN(n510) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n507) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT104), .B(n508), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n511), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n561), .A2(n521), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n521), .ZN(n516) );
  XOR2_X1 U580 ( .A(KEYINPUT108), .B(n516), .Z(n517) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n527), .A2(n521), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n523) );
  NOR2_X1 U587 ( .A1(n529), .A2(n521), .ZN(n522) );
  XOR2_X1 U588 ( .A(n523), .B(n522), .Z(G1339GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n561), .ZN(n525) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n541) );
  NOR2_X1 U591 ( .A1(n527), .A2(n541), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT114), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT115), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n564), .A2(n537), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U598 ( .A1(n537), .A2(n545), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n557), .A2(n537), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NAND2_X1 U603 ( .A1(n537), .A2(n552), .ZN(n539) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n538) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n544) );
  NOR2_X1 U607 ( .A1(n559), .A2(n541), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(n542), .Z(n551) );
  NAND2_X1 U609 ( .A1(n564), .A2(n551), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  NAND2_X1 U612 ( .A1(n551), .A2(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n343), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n564), .A2(n556), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n555), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  INV_X1 U626 ( .A(n559), .ZN(n560) );
  AND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  AND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n574), .A2(n564), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U633 ( .A1(n574), .A2(n568), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(n571), .ZN(G1353GAT) );
  XOR2_X1 U636 ( .A(G211GAT), .B(KEYINPUT127), .Z(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n343), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  INV_X1 U639 ( .A(n574), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

