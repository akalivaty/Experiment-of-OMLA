

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X2 U323 ( .A(n461), .B(n438), .ZN(n567) );
  XNOR2_X1 U324 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U325 ( .A(n474), .B(KEYINPUT118), .ZN(n475) );
  XNOR2_X1 U326 ( .A(n368), .B(n367), .ZN(n580) );
  XNOR2_X1 U327 ( .A(n366), .B(KEYINPUT89), .ZN(n367) );
  XNOR2_X1 U328 ( .A(n436), .B(n355), .ZN(n356) );
  XNOR2_X1 U329 ( .A(n422), .B(KEYINPUT37), .ZN(n490) );
  XNOR2_X1 U330 ( .A(n363), .B(n362), .ZN(n541) );
  XNOR2_X1 U331 ( .A(n343), .B(n342), .ZN(n352) );
  XNOR2_X1 U332 ( .A(n444), .B(n292), .ZN(n342) );
  XOR2_X1 U333 ( .A(KEYINPUT47), .B(n468), .Z(n291) );
  AND2_X1 U334 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U335 ( .A(G15GAT), .B(n353), .Z(n293) );
  INV_X1 U336 ( .A(G183GAT), .ZN(n385) );
  XNOR2_X1 U337 ( .A(n386), .B(n385), .ZN(n387) );
  INV_X1 U338 ( .A(KEYINPUT108), .ZN(n470) );
  INV_X1 U339 ( .A(KEYINPUT92), .ZN(n374) );
  XNOR2_X1 U340 ( .A(n431), .B(n387), .ZN(n388) );
  XNOR2_X1 U341 ( .A(n470), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U342 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U343 ( .A(n472), .B(n471), .ZN(n538) );
  XNOR2_X1 U344 ( .A(n398), .B(n397), .ZN(n401) );
  INV_X1 U345 ( .A(n490), .ZN(n491) );
  XNOR2_X1 U346 ( .A(n357), .B(n356), .ZN(n363) );
  XOR2_X1 U347 ( .A(n403), .B(n402), .Z(n589) );
  INV_X1 U348 ( .A(G190GAT), .ZN(n485) );
  XNOR2_X1 U349 ( .A(n493), .B(n492), .ZN(n513) );
  XNOR2_X1 U350 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U351 ( .A(n456), .B(G106GAT), .ZN(n457) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U353 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U354 ( .A(n495), .B(n494), .ZN(G1330GAT) );
  XOR2_X1 U355 ( .A(KEYINPUT82), .B(KEYINPUT86), .Z(n295) );
  XNOR2_X1 U356 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U358 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n297) );
  XNOR2_X1 U359 ( .A(KEYINPUT5), .B(G1GAT), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U361 ( .A(n299), .B(n298), .Z(n305) );
  XNOR2_X1 U362 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n300), .B(KEYINPUT2), .ZN(n318) );
  XOR2_X1 U364 ( .A(G162GAT), .B(n318), .Z(n302) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U366 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G148GAT), .Z(n307) );
  XNOR2_X1 U370 ( .A(G85GAT), .B(G120GAT), .ZN(n306) );
  XNOR2_X1 U371 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U372 ( .A(n309), .B(n308), .Z(n317) );
  XOR2_X1 U373 ( .A(KEYINPUT0), .B(G134GAT), .Z(n311) );
  XNOR2_X1 U374 ( .A(G127GAT), .B(G113GAT), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U376 ( .A(KEYINPUT78), .B(n312), .Z(n361) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT1), .Z(n314) );
  XNOR2_X1 U378 ( .A(KEYINPUT83), .B(KEYINPUT6), .ZN(n313) );
  XNOR2_X1 U379 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U380 ( .A(n361), .B(n315), .ZN(n316) );
  XNOR2_X1 U381 ( .A(n317), .B(n316), .ZN(n529) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G50GAT), .Z(n417) );
  XNOR2_X1 U383 ( .A(n417), .B(n318), .ZN(n320) );
  AND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n321), .B(KEYINPUT22), .ZN(n323) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G22GAT), .Z(n442) );
  XOR2_X1 U388 ( .A(G218GAT), .B(n442), .Z(n322) );
  XNOR2_X1 U389 ( .A(n323), .B(n322), .ZN(n333) );
  XOR2_X1 U390 ( .A(G197GAT), .B(KEYINPUT21), .Z(n325) );
  XNOR2_X1 U391 ( .A(G211GAT), .B(KEYINPUT80), .ZN(n324) );
  XNOR2_X1 U392 ( .A(n325), .B(n324), .ZN(n350) );
  INV_X1 U393 ( .A(G78GAT), .ZN(n326) );
  NAND2_X1 U394 ( .A1(G204GAT), .A2(n326), .ZN(n329) );
  INV_X1 U395 ( .A(G204GAT), .ZN(n327) );
  NAND2_X1 U396 ( .A1(n327), .A2(G78GAT), .ZN(n328) );
  NAND2_X1 U397 ( .A1(n329), .A2(n328), .ZN(n331) );
  XNOR2_X1 U398 ( .A(G148GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U399 ( .A(n331), .B(n330), .ZN(n423) );
  XNOR2_X1 U400 ( .A(n350), .B(n423), .ZN(n332) );
  XNOR2_X1 U401 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U402 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n335) );
  XNOR2_X1 U403 ( .A(KEYINPUT79), .B(KEYINPUT81), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n478) );
  XOR2_X1 U406 ( .A(KEYINPUT88), .B(G204GAT), .Z(n341) );
  XNOR2_X1 U407 ( .A(G218GAT), .B(G36GAT), .ZN(n338) );
  XNOR2_X1 U408 ( .A(n338), .B(G190GAT), .ZN(n410) );
  XNOR2_X1 U409 ( .A(G92GAT), .B(G64GAT), .ZN(n339) );
  XNOR2_X1 U410 ( .A(n339), .B(G176GAT), .ZN(n430) );
  XNOR2_X1 U411 ( .A(n410), .B(n430), .ZN(n340) );
  XNOR2_X1 U412 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G169GAT), .Z(n444) );
  INV_X1 U414 ( .A(KEYINPUT17), .ZN(n344) );
  NAND2_X1 U415 ( .A1(KEYINPUT18), .A2(n344), .ZN(n347) );
  INV_X1 U416 ( .A(KEYINPUT18), .ZN(n345) );
  NAND2_X1 U417 ( .A1(n345), .A2(KEYINPUT17), .ZN(n346) );
  NAND2_X1 U418 ( .A1(n347), .A2(n346), .ZN(n349) );
  XNOR2_X1 U419 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n348) );
  XNOR2_X1 U420 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U421 ( .A(n353), .B(n350), .Z(n351) );
  XNOR2_X1 U422 ( .A(n352), .B(n351), .ZN(n533) );
  NAND2_X1 U423 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U424 ( .A(n293), .B(n354), .ZN(n357) );
  XNOR2_X1 U425 ( .A(G120GAT), .B(G71GAT), .ZN(n436) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(G190GAT), .ZN(n355) );
  XOR2_X1 U427 ( .A(G176GAT), .B(KEYINPUT20), .Z(n359) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(G169GAT), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U431 ( .A1(n533), .A2(n541), .ZN(n364) );
  NAND2_X1 U432 ( .A1(n478), .A2(n364), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n365), .B(KEYINPUT25), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n533), .B(KEYINPUT27), .ZN(n377) );
  INV_X1 U435 ( .A(n377), .ZN(n369) );
  OR2_X1 U436 ( .A1(n478), .A2(n541), .ZN(n368) );
  XOR2_X1 U437 ( .A(KEYINPUT90), .B(KEYINPUT26), .Z(n366) );
  NOR2_X1 U438 ( .A1(n369), .A2(n580), .ZN(n370) );
  NOR2_X1 U439 ( .A1(n371), .A2(n370), .ZN(n372) );
  XOR2_X1 U440 ( .A(KEYINPUT91), .B(n372), .Z(n373) );
  NOR2_X1 U441 ( .A1(n529), .A2(n373), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U443 ( .A(n478), .B(KEYINPUT65), .Z(n376) );
  XNOR2_X1 U444 ( .A(n376), .B(KEYINPUT28), .ZN(n540) );
  NAND2_X1 U445 ( .A1(n529), .A2(n377), .ZN(n537) );
  NOR2_X1 U446 ( .A1(n537), .A2(n541), .ZN(n378) );
  NAND2_X1 U447 ( .A1(n540), .A2(n378), .ZN(n379) );
  NAND2_X1 U448 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n381), .B(KEYINPUT93), .ZN(n498) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n383) );
  XNOR2_X1 U451 ( .A(KEYINPUT76), .B(KEYINPUT74), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n383), .B(n382), .ZN(n403) );
  XNOR2_X1 U453 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n384), .B(KEYINPUT70), .ZN(n431) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(G71GAT), .B(n388), .ZN(n398) );
  XOR2_X1 U457 ( .A(G22GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U458 ( .A(G127GAT), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U460 ( .A(G8GAT), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT75), .ZN(n391) );
  XNOR2_X1 U462 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U463 ( .A(n394), .B(n393), .Z(n396) );
  INV_X1 U464 ( .A(KEYINPUT15), .ZN(n395) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(G15GAT), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n399), .B(KEYINPUT68), .ZN(n445) );
  XNOR2_X1 U467 ( .A(n445), .B(KEYINPUT14), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U469 ( .A1(n498), .A2(n589), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n404), .B(KEYINPUT96), .ZN(n420) );
  XOR2_X1 U471 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n406) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U474 ( .A(n407), .B(KEYINPUT9), .Z(n412) );
  XOR2_X1 U475 ( .A(G43GAT), .B(KEYINPUT7), .Z(n409) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n439) );
  XNOR2_X1 U478 ( .A(n439), .B(n410), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U480 ( .A(G92GAT), .B(G106GAT), .Z(n414) );
  XNOR2_X1 U481 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U483 ( .A(n416), .B(n415), .Z(n419) );
  XOR2_X1 U484 ( .A(G85GAT), .B(G99GAT), .Z(n435) );
  XNOR2_X1 U485 ( .A(n417), .B(n435), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n564) );
  XNOR2_X1 U487 ( .A(KEYINPUT36), .B(n564), .ZN(n593) );
  NAND2_X1 U488 ( .A1(n420), .A2(n593), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n421), .B(KEYINPUT97), .ZN(n422) );
  XOR2_X1 U490 ( .A(n423), .B(KEYINPUT72), .Z(n425) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U493 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n427) );
  XNOR2_X1 U494 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U496 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n461) );
  XOR2_X1 U501 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n438) );
  XOR2_X1 U502 ( .A(n439), .B(KEYINPUT69), .Z(n441) );
  NAND2_X1 U503 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U505 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n455) );
  XOR2_X1 U508 ( .A(G197GAT), .B(G36GAT), .Z(n449) );
  XNOR2_X1 U509 ( .A(G113GAT), .B(G50GAT), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n451) );
  XNOR2_X1 U512 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U514 ( .A(n453), .B(n452), .Z(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n489) );
  NAND2_X1 U516 ( .A1(n567), .A2(n489), .ZN(n518) );
  NOR2_X1 U517 ( .A1(n490), .A2(n518), .ZN(n535) );
  INV_X1 U518 ( .A(n540), .ZN(n524) );
  NAND2_X1 U519 ( .A1(n535), .A2(n524), .ZN(n458) );
  XOR2_X1 U520 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n456) );
  XNOR2_X1 U521 ( .A(n458), .B(n457), .ZN(G1339GAT) );
  XOR2_X1 U522 ( .A(KEYINPUT45), .B(KEYINPUT107), .Z(n460) );
  NAND2_X1 U523 ( .A1(n589), .A2(n593), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n460), .B(n459), .ZN(n462) );
  NOR2_X1 U525 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n489), .A2(n463), .ZN(n469) );
  INV_X1 U527 ( .A(n489), .ZN(n581) );
  NAND2_X1 U528 ( .A1(n581), .A2(n567), .ZN(n464) );
  XNOR2_X1 U529 ( .A(KEYINPUT46), .B(n464), .ZN(n466) );
  NOR2_X1 U530 ( .A1(n564), .A2(n589), .ZN(n465) );
  NAND2_X1 U531 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U532 ( .A(KEYINPUT106), .B(n467), .ZN(n468) );
  NAND2_X1 U533 ( .A1(n469), .A2(n291), .ZN(n472) );
  INV_X1 U534 ( .A(n538), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n473), .A2(n533), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n474) );
  NOR2_X1 U537 ( .A1(n477), .A2(n529), .ZN(n578) );
  NAND2_X1 U538 ( .A1(n578), .A2(n478), .ZN(n479) );
  XNOR2_X1 U539 ( .A(KEYINPUT55), .B(n479), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n480), .A2(n541), .ZN(n574) );
  NOR2_X1 U541 ( .A1(n489), .A2(n574), .ZN(n483) );
  XNOR2_X1 U542 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n481), .B(G169GAT), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1348GAT) );
  INV_X1 U545 ( .A(n564), .ZN(n484) );
  NOR2_X1 U546 ( .A1(n574), .A2(n484), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n486) );
  NOR2_X1 U548 ( .A1(n489), .A2(n461), .ZN(n499) );
  NAND2_X1 U549 ( .A1(n499), .A2(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n492) );
  NAND2_X1 U551 ( .A1(n513), .A2(n541), .ZN(n495) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n501) );
  INV_X1 U553 ( .A(n589), .ZN(n575) );
  NOR2_X1 U554 ( .A1(n564), .A2(n575), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  NOR2_X1 U556 ( .A1(n498), .A2(n497), .ZN(n516) );
  AND2_X1 U557 ( .A1(n499), .A2(n516), .ZN(n506) );
  NAND2_X1 U558 ( .A1(n506), .A2(n529), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U560 ( .A(G1GAT), .B(n502), .Z(G1324GAT) );
  NAND2_X1 U561 ( .A1(n533), .A2(n506), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U564 ( .A1(n506), .A2(n541), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U566 ( .A1(n524), .A2(n506), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U568 ( .A1(n513), .A2(n529), .ZN(n510) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(KEYINPUT95), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  XOR2_X1 U572 ( .A(G36GAT), .B(KEYINPUT99), .Z(n512) );
  NAND2_X1 U573 ( .A1(n513), .A2(n533), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1329GAT) );
  XNOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT100), .ZN(n515) );
  NAND2_X1 U576 ( .A1(n513), .A2(n524), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n520) );
  INV_X1 U579 ( .A(n516), .ZN(n517) );
  NOR2_X1 U580 ( .A1(n518), .A2(n517), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n525), .A2(n529), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U584 ( .A1(n533), .A2(n525), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n541), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U592 ( .A1(n535), .A2(n529), .ZN(n532) );
  XOR2_X1 U593 ( .A(G85GAT), .B(KEYINPUT103), .Z(n530) );
  XNOR2_X1 U594 ( .A(KEYINPUT104), .B(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n535), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n535), .A2(n541), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT109), .B(n539), .ZN(n554) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n554), .A2(n542), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n549), .A2(n581), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT110), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U608 ( .A1(n549), .A2(n567), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n549), .A2(n589), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT111), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U614 ( .A1(n549), .A2(n564), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT112), .Z(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NOR2_X1 U618 ( .A1(n580), .A2(n554), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT113), .B(n555), .Z(n565) );
  NAND2_X1 U620 ( .A1(n581), .A2(n565), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT114), .B(n559), .Z(n561) );
  NAND2_X1 U626 ( .A1(n565), .A2(n567), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n589), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT116), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U633 ( .A(n567), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n568), .A2(n574), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT121), .B(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1350GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n592) );
  AND2_X1 U645 ( .A1(n581), .A2(n592), .ZN(n583) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U651 ( .A1(n592), .A2(n461), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G204GAT), .ZN(G1353GAT) );
  XOR2_X1 U654 ( .A(G211GAT), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1354GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT62), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

