//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n461), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT67), .ZN(G160));
  NOR2_X1   g050(.A1(new_n464), .A2(new_n469), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n476), .B(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(new_n465), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n465), .A2(KEYINPUT68), .A3(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n470), .A2(KEYINPUT71), .A3(G138), .A4(new_n469), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(KEYINPUT71), .A3(KEYINPUT4), .A4(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n469), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n476), .A2(G126), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n492), .A2(new_n493), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .A3(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT73), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n511), .A2(new_n514), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n510), .A2(G51), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT74), .B(G89), .Z(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(new_n526), .B1(new_n512), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n513), .A2(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n510), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT5), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n531), .A2(new_n532), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND4_X1  g118(.A1(new_n508), .A2(G43), .A3(G543), .A4(new_n509), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n508), .A2(new_n509), .A3(new_n512), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(KEYINPUT75), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n504), .B1(new_n548), .B2(KEYINPUT75), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n508), .A2(G543), .A3(new_n509), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n562), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n508), .A2(G91), .A3(new_n509), .A4(new_n512), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n567), .B2(new_n504), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n510), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n562), .A2(G87), .A3(new_n512), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n510), .A2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n513), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n538), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n538), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n510), .A2(G47), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n513), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(KEYINPUT76), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n559), .A2(new_n594), .B1(new_n595), .B2(new_n504), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n508), .A2(G92), .A3(new_n509), .A4(new_n512), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n562), .A2(KEYINPUT10), .A3(G92), .A4(new_n512), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n568), .B1(new_n561), .B2(new_n564), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(G868), .B2(new_n605), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(G868), .B2(new_n605), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n513), .A2(G81), .ZN(new_n610));
  NAND2_X1  g185(.A1(G68), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G56), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n538), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n610), .B(new_n544), .C1(new_n615), .C2(new_n549), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n599), .A2(new_n600), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n535), .A2(new_n537), .A3(G66), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n504), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n510), .B2(G54), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(new_n617), .ZN(G323));
  XOR2_X1   g201(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n627));
  XNOR2_X1  g202(.A(G323), .B(new_n627), .ZN(G282));
  NAND2_X1  g203(.A1(new_n470), .A2(new_n466), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n631), .A2(new_n632), .B1(KEYINPUT78), .B2(G2100), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  OR3_X1    g209(.A1(new_n634), .A2(KEYINPUT78), .A3(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n481), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n478), .B2(G123), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(KEYINPUT78), .B2(G2100), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n641), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  INV_X1    g219(.A(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT79), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT16), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n650), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2443), .B(G2446), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n658), .A3(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n662), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n668), .A2(new_n669), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT81), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT82), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n686), .A2(KEYINPUT82), .A3(new_n692), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n691), .B(new_n693), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1991), .ZN(new_n698));
  INV_X1    g273(.A(G1996), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n697), .A2(G1991), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(G1991), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(G1996), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n702), .B1(new_n700), .B2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n683), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n710), .A2(new_n682), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(G229));
  NAND2_X1  g287(.A1(new_n640), .A2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT30), .B(G28), .Z(new_n714));
  NOR2_X1   g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n713), .B1(G29), .B2(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  NOR2_X1   g293(.A1(G5), .A2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G171), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G35), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT93), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(G2090), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT23), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT84), .B(G16), .ZN(new_n732));
  INV_X1    g307(.A(G20), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n731), .B(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G16), .B2(G299), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1956), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n728), .A2(KEYINPUT94), .A3(G2090), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n727), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n729), .B(new_n737), .C1(new_n738), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G160), .A2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G34), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n745), .B1(G29), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n751), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n465), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n466), .A2(G105), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n478), .B2(G129), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G27), .A2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G164), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n601), .B2(G16), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n765), .B(new_n769), .C1(G1348), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n748), .A2(new_n749), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n753), .A2(G1966), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n755), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n776), .A2(G29), .A3(G33), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(G29), .B2(G33), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n469), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n466), .A2(G103), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n465), .A2(G139), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n783), .A2(KEYINPUT89), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(KEYINPUT89), .B1(new_n783), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n777), .B(new_n778), .C1(new_n791), .C2(new_n724), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2072), .ZN(new_n793));
  INV_X1    g368(.A(G19), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n732), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n616), .B2(new_n732), .ZN(new_n796));
  INV_X1    g371(.A(G1341), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n771), .A2(G1348), .ZN(new_n799));
  AOI21_X1  g374(.A(KEYINPUT28), .B1(new_n724), .B2(G26), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n724), .A2(G26), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n465), .A2(G140), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n469), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n478), .B2(G128), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n801), .B1(new_n806), .B2(new_n724), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(KEYINPUT28), .ZN(new_n808));
  INV_X1    g383(.A(G2067), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n799), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI211_X1 g385(.A(new_n798), .B(new_n810), .C1(new_n809), .C2(new_n808), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n775), .A2(new_n793), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n744), .A2(new_n812), .ZN(new_n813));
  MUX2_X1   g388(.A(G22), .B(G303), .S(new_n732), .Z(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G1971), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n751), .A2(G6), .ZN(new_n816));
  INV_X1    g391(.A(G305), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n751), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT32), .B(G1981), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G16), .A2(G23), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT86), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G288), .B2(new_n751), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT33), .B(G1976), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n815), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT34), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n732), .A2(G24), .ZN(new_n829));
  XNOR2_X1  g404(.A(G290), .B(KEYINPUT85), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n732), .ZN(new_n831));
  INV_X1    g406(.A(G1986), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n724), .A2(G25), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n465), .A2(G131), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n469), .A2(G107), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n478), .B2(G119), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n834), .B1(new_n839), .B2(new_n724), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G1991), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT83), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(KEYINPUT87), .B2(KEYINPUT36), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n828), .A2(new_n833), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n828), .A2(new_n848), .A3(new_n833), .A4(new_n844), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n813), .A2(new_n847), .A3(new_n849), .ZN(G150));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g426(.A1(G150), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n813), .A2(new_n847), .A3(KEYINPUT97), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(G311));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n535), .A2(new_n537), .A3(G67), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n856), .A2(KEYINPUT99), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT99), .B1(new_n856), .B2(new_n857), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n508), .A2(G55), .A3(G543), .A4(new_n509), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n508), .A2(G93), .A3(new_n509), .A4(new_n512), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n855), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n856), .A2(new_n857), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(G651), .A3(new_n858), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n862), .A2(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G860), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT102), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n552), .B1(new_n865), .B2(new_n871), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n616), .B1(new_n869), .B2(new_n870), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT101), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT100), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT100), .B1(new_n869), .B2(new_n870), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n616), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n624), .A2(new_n608), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT39), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n887), .B(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(G860), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n886), .A2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n876), .B1(new_n892), .B2(new_n893), .ZN(G145));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n787), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n478), .A2(G129), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n806), .B1(new_n897), .B2(new_n761), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n478), .A2(G128), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n762), .B1(new_n899), .B2(new_n805), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n900), .A3(G164), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G164), .B1(new_n900), .B2(new_n898), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n791), .B(new_n896), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n901), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n904), .B2(new_n907), .ZN(new_n911));
  OAI21_X1  g486(.A(G162), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n631), .B(new_n839), .ZN(new_n913));
  XNOR2_X1  g488(.A(G160), .B(new_n640), .ZN(new_n914));
  OR2_X1    g489(.A1(G106), .A2(G2105), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n915), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n916));
  INV_X1    g491(.A(G142), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n481), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n478), .B2(G130), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n914), .A2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  INV_X1    g499(.A(new_n913), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n904), .A2(new_n907), .ZN(new_n928));
  INV_X1    g503(.A(new_n908), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n909), .A3(new_n488), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n912), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n912), .B2(new_n931), .ZN(new_n935));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n936));
  OR3_X1    g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G395));
  XOR2_X1   g514(.A(new_n885), .B(new_n625), .Z(new_n940));
  NAND2_X1  g515(.A1(new_n601), .A2(G299), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n605), .A2(new_n624), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT41), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n601), .A2(G299), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n605), .A2(new_n624), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n941), .A2(new_n942), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT107), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n940), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT42), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G290), .A2(new_n574), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n590), .A2(G288), .A3(new_n591), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT110), .ZN(new_n960));
  XNOR2_X1  g535(.A(G303), .B(KEYINPUT109), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(new_n817), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n963), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n961), .B(G305), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n959), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n950), .B(new_n970), .C1(new_n940), .C2(new_n954), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n956), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n956), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(G868), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n873), .A2(new_n617), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n975), .ZN(G331));
  XOR2_X1   g552(.A(G286), .B(G301), .Z(new_n978));
  OAI21_X1  g553(.A(new_n552), .B1(new_n861), .B2(new_n864), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n883), .B1(new_n882), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G286), .B(G301), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n879), .A2(new_n884), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n982), .A2(new_n952), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n948), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n980), .A2(new_n981), .A3(new_n978), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n879), .B2(new_n884), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n949), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n969), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n947), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n944), .B2(new_n945), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n952), .A2(KEYINPUT113), .A3(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1000), .B(new_n1001), .C1(new_n988), .C2(new_n989), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n982), .A2(new_n953), .A3(new_n984), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n982), .A2(new_n984), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1001), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n968), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n993), .A2(new_n1007), .A3(new_n933), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n982), .A2(new_n952), .A3(new_n984), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n991), .B1(new_n990), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n986), .A2(KEYINPUT112), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n968), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n993), .A3(new_n1016), .A4(new_n933), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1017), .A2(KEYINPUT44), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(KEYINPUT115), .A3(KEYINPUT43), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1011), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1022));
  AOI21_X1  g597(.A(G37), .B1(new_n1022), .B2(new_n969), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1016), .B1(new_n1023), .B2(new_n1015), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1020), .A2(new_n1026), .ZN(G397));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n471), .A2(new_n472), .ZN(new_n1031));
  OAI211_X1 g606(.A(G40), .B(new_n467), .C1(new_n1031), .C2(new_n469), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n806), .B(G2067), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n762), .B(G1996), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n842), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n839), .B(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G290), .A2(G1986), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n832), .B1(new_n590), .B2(new_n591), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1033), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n501), .A2(new_n1028), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n468), .A2(new_n473), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1045), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G305), .A2(G1981), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT117), .B(G1981), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n576), .A2(new_n577), .A3(new_n581), .A4(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n573), .A2(new_n572), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n571), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1055), .A2(new_n571), .A3(KEYINPUT118), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1051), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1054), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1053), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1049), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G303), .A2(G8), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n501), .A2(new_n1028), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT50), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n501), .A2(new_n1071), .A3(new_n1028), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n742), .A2(new_n1070), .A3(new_n1048), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT45), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1032), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1028), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1971), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1068), .B(G8), .C1(new_n1073), .C2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1048), .A2(new_n1028), .A3(new_n501), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n574), .A2(new_n1080), .A3(G1976), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1055), .A2(G1976), .A3(new_n571), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT116), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .A4(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT52), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1049), .A2(new_n1081), .A3(new_n1086), .A4(new_n1083), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1049), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1065), .B1(new_n1078), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT119), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1065), .B(new_n1092), .C1(new_n1078), .C2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1028), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1095), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1070), .A2(new_n1048), .A3(new_n1072), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1096), .A2(G1966), .B1(new_n1097), .B2(G2084), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(G8), .A3(G168), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1089), .B1(new_n1099), .B2(KEYINPUT121), .ZN(new_n1100));
  OAI21_X1  g675(.A(G8), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1067), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1098), .A2(new_n1103), .A3(G8), .A4(G168), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(new_n1102), .A3(new_n1078), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1094), .B1(KEYINPUT63), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1078), .A2(KEYINPUT120), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1096), .A2(G1971), .B1(new_n1097), .B2(G2090), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1068), .B1(new_n1108), .B2(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(KEYINPUT120), .A3(new_n1078), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT63), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1104), .A3(new_n1100), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G299), .B(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1097), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1075), .A2(new_n1076), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1114), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1097), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G1348), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1048), .A2(new_n1028), .A3(new_n809), .A4(new_n501), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT122), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n601), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1117), .A2(new_n1119), .A3(new_n1114), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1120), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1123), .B(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1129), .C1(G1348), .C2(new_n1121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1128), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1096), .A2(new_n699), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(new_n797), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1079), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1079), .A2(KEYINPUT124), .A3(new_n1138), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1143), .A2(KEYINPUT59), .A3(new_n552), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT59), .B1(new_n1143), .B2(new_n552), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1135), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1114), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1119), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1116), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT61), .B1(new_n1126), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1147), .A3(new_n1116), .ZN(new_n1151));
  NOR2_X1   g726(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1120), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1149), .A2(KEYINPUT125), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1127), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1089), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1075), .A2(new_n768), .A3(new_n1076), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1097), .A2(new_n721), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n768), .A4(new_n1076), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1160), .A2(new_n1161), .A3(G301), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT54), .B1(new_n1164), .B2(KEYINPUT126), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1162), .A3(new_n1161), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(new_n1163), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G168), .A2(new_n1045), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AND4_X1   g747(.A1(new_n749), .A2(new_n1070), .A3(new_n1048), .A4(new_n1072), .ZN(new_n1173));
  AOI21_X1  g748(.A(G1966), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT51), .B(new_n1172), .C1(new_n1175), .C2(new_n1045), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1098), .A2(new_n1171), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT51), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1178), .B(G8), .C1(new_n1098), .C2(G286), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1167), .A2(KEYINPUT54), .A3(new_n1163), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1157), .A2(new_n1170), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1106), .B(new_n1113), .C1(new_n1156), .C2(new_n1182), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1180), .A2(KEYINPUT62), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1089), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1186));
  AOI211_X1 g761(.A(KEYINPUT120), .B(new_n1068), .C1(new_n1108), .C2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1176), .A2(new_n1179), .A3(new_n1189), .A4(new_n1177), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1167), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT127), .B1(new_n1188), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1157), .A2(new_n1194), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1184), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1044), .B1(new_n1183), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1033), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1198), .B1(new_n1034), .B2(new_n762), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1033), .A2(new_n699), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT47), .Z(new_n1204));
  AND4_X1   g779(.A1(new_n1037), .A2(new_n1034), .A3(new_n1035), .A4(new_n839), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1205), .B1(new_n809), .B2(new_n806), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1198), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1041), .A2(new_n1198), .ZN(new_n1208));
  OR2_X1    g783(.A1(new_n1208), .A2(KEYINPUT48), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(new_n1198), .B2(new_n1039), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1210), .B1(KEYINPUT48), .B2(new_n1208), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1204), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1197), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g788(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1215));
  NOR2_X1   g789(.A1(G227), .A2(new_n458), .ZN(new_n1216));
  AND4_X1   g790(.A1(new_n666), .A2(new_n709), .A3(new_n711), .A4(new_n1216), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1217), .B1(new_n934), .B2(new_n935), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1215), .A2(new_n1218), .ZN(G308));
  OAI221_X1 g793(.A(new_n1217), .B1(new_n934), .B2(new_n935), .C1(new_n1024), .C2(new_n1025), .ZN(G225));
endmodule


