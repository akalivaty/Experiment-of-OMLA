//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT66), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT67), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT70), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G169), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G283), .ZN(new_n251));
  INV_X1    g0051(.A(G97), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n251), .B(new_n207), .C1(G33), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n213), .ZN(new_n255));
  INV_X1    g0055(.A(G116), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT20), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n207), .A3(G1), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G116), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n262), .A2(new_n255), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n267), .B2(G116), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n250), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  OAI211_X1 g0073(.A(G257), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n265), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n272), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n206), .A2(G45), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT5), .A2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT5), .A2(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n213), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n280), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT5), .B(G41), .ZN(new_n293));
  INV_X1    g0093(.A(new_n285), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n281), .ZN(new_n296));
  INV_X1    g0096(.A(G270), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT84), .B1(new_n284), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n293), .A2(new_n294), .B1(new_n290), .B2(new_n280), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G270), .B1(new_n288), .B2(new_n291), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT84), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n283), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n269), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT21), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n301), .A2(new_n302), .A3(new_n283), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n302), .B1(new_n301), .B2(new_n283), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT21), .A3(new_n269), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n260), .A2(new_n268), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n301), .A2(G179), .A3(new_n283), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n306), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G190), .B1(new_n307), .B2(new_n308), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n299), .A2(G200), .A3(new_n303), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n311), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(KEYINPUT85), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT85), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n306), .A2(new_n310), .A3(new_n314), .ZN(new_n321));
  INV_X1    g0121(.A(new_n318), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n203), .A2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G20), .A2(G33), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n265), .A2(G20), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n325), .B1(new_n326), .B2(new_n328), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n255), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n262), .A2(new_n255), .ZN(new_n334));
  INV_X1    g0134(.A(G50), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n206), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n334), .A2(new_n336), .B1(new_n335), .B2(new_n262), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT9), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n281), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT72), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT72), .B1(new_n281), .B2(new_n340), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT71), .B(G226), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n276), .A2(new_n277), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G222), .A3(new_n273), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G223), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n349), .B1(new_n350), .B2(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n282), .ZN(new_n354));
  INV_X1    g0154(.A(new_n340), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n281), .A3(G274), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n347), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(G200), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n339), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n339), .A2(new_n363), .A3(new_n359), .A4(new_n360), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n357), .A2(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT73), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n357), .B2(new_n250), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n367), .B(new_n338), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n262), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n327), .A2(G50), .B1(G20), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n330), .B2(new_n350), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n206), .A2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n334), .A2(G68), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT11), .B1(new_n376), .B2(new_n255), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n348), .A2(G226), .A3(new_n273), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n348), .A2(KEYINPUT74), .A3(G226), .A4(new_n273), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT76), .B1(new_n265), .B2(new_n252), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(G33), .A3(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n348), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n388), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n282), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g0200(.A(G238), .B1(new_n343), .B2(new_n344), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n356), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n281), .B1(new_n388), .B2(new_n397), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT13), .B1(new_n405), .B2(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G169), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(G179), .A3(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n407), .B2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n383), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n382), .B1(new_n407), .B2(new_n358), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n404), .B2(new_n406), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n345), .A2(G244), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n348), .A2(G232), .A3(new_n273), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  INV_X1    g0222(.A(G238), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n421), .B1(new_n422), .B2(new_n348), .C1(new_n351), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n282), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n425), .A3(new_n356), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n331), .A2(new_n328), .B1(new_n207), .B2(new_n350), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT15), .B(G87), .Z(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n329), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n255), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n334), .A2(G77), .A3(new_n378), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G77), .B2(new_n263), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n426), .B2(new_n250), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n427), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n426), .A2(G200), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n435), .B1(new_n426), .B2(new_n358), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n371), .A2(new_n419), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n331), .B1(new_n206), .B2(G20), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n334), .B1(new_n262), .B2(new_n331), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n352), .A2(new_n273), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n444), .B1(G226), .B2(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G87), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n281), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G232), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n356), .B1(new_n341), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n415), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n447), .A2(new_n450), .A3(new_n358), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(G58), .A2(G68), .ZN(new_n455));
  OAI21_X1  g0255(.A(G20), .B1(new_n455), .B2(new_n202), .ZN(new_n456));
  INV_X1    g0256(.A(G159), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n457), .A2(KEYINPUT78), .A3(G20), .A4(G33), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT78), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n327), .B2(G159), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT16), .B(new_n456), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n270), .A2(new_n271), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(new_n207), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n276), .A2(new_n207), .A3(new_n277), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT7), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n469), .A3(G68), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n431), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT16), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n466), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n277), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n372), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n471), .B2(new_n477), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n443), .B(new_n454), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT17), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n481), .B(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n443), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n447), .A2(new_n450), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G179), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n250), .B2(new_n485), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(KEYINPUT18), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT18), .ZN(new_n491));
  INV_X1    g0291(.A(new_n443), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n462), .A2(new_n470), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n255), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n270), .A2(new_n271), .A3(G20), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n474), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G68), .ZN(new_n498));
  INV_X1    g0298(.A(new_n476), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT16), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT79), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n492), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n487), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n491), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n484), .A2(KEYINPUT80), .A3(KEYINPUT18), .A4(new_n487), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n490), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n490), .A2(KEYINPUT81), .A3(new_n505), .A4(new_n506), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n483), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n441), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n348), .A2(G257), .A3(G1698), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G294), .ZN(new_n515));
  OAI211_X1 g0315(.A(G250), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n282), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n300), .A2(G264), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n292), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n415), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n518), .A2(new_n358), .A3(new_n292), .A4(new_n519), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT25), .B1(new_n262), .B2(new_n422), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n422), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(new_n267), .B2(G107), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n207), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n528));
  AND2_X1   g0328(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n348), .A2(new_n207), .A3(G87), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n207), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n422), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n532), .A2(new_n533), .A3(new_n542), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT87), .B1(new_n544), .B2(new_n255), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n546), .B(new_n431), .C1(new_n541), .C2(new_n543), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n523), .B(new_n527), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n527), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n255), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n546), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n255), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n520), .A2(new_n250), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(G179), .B2(new_n520), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n548), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT88), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n527), .B1(new_n545), .B2(new_n547), .ZN(new_n558));
  INV_X1    g0358(.A(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT88), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n548), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n263), .A2(G97), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n267), .B2(G97), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT6), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n567), .A2(new_n252), .A3(G107), .ZN(new_n568));
  XNOR2_X1  g0368(.A(G97), .B(G107), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(new_n207), .B1(new_n350), .B2(new_n328), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n422), .B1(new_n473), .B2(new_n474), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n255), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT82), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n255), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n566), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n295), .A2(G257), .A3(new_n281), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n292), .ZN(new_n580));
  OAI211_X1 g0380(.A(G244), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n348), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n348), .A2(G250), .A3(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n251), .A4(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n580), .B1(new_n282), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G169), .ZN(new_n588));
  INV_X1    g0388(.A(G179), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n587), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n578), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(G190), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n577), .B(new_n592), .C1(new_n415), .C2(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT19), .B1(new_n329), .B2(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n463), .A2(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(G68), .ZN(new_n597));
  INV_X1    g0397(.A(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(new_n252), .A3(new_n422), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT19), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n389), .B2(new_n391), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n601), .B2(G20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n429), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n255), .B1(new_n262), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n267), .A2(new_n429), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n607));
  OAI211_X1 g0407(.A(G238), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n534), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n282), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n294), .A2(new_n281), .A3(G274), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n281), .A2(G250), .A3(new_n285), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT83), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n610), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n605), .A2(new_n606), .B1(new_n617), .B2(new_n589), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n614), .A3(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n250), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(G200), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n267), .A2(G87), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n610), .A2(new_n614), .A3(G190), .A4(new_n616), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n605), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n594), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n324), .A2(new_n513), .A3(new_n563), .A4(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n437), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n418), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n483), .B1(new_n630), .B2(new_n413), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n505), .A2(new_n488), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n365), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(new_n370), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n605), .A2(new_n623), .A3(new_n624), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n609), .A2(new_n636), .A3(new_n282), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n609), .B2(new_n282), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n616), .B(new_n614), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n250), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n635), .A2(new_n640), .B1(new_n618), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n591), .A2(new_n642), .A3(new_n593), .A4(new_n548), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n321), .B1(new_n558), .B2(new_n559), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n578), .A2(new_n621), .A3(new_n590), .A4(new_n625), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT26), .ZN(new_n647));
  INV_X1    g0447(.A(new_n587), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(G179), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n577), .A2(new_n649), .A3(new_n588), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n618), .A2(new_n641), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n634), .B1(new_n512), .B2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n563), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n553), .A2(new_n664), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n657), .A2(new_n665), .B1(new_n560), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n324), .B1(new_n311), .B2(new_n664), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n321), .A2(new_n312), .A3(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n669), .A3(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n315), .A2(new_n663), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n563), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n558), .A2(new_n559), .A3(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n210), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n599), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n681), .A2(KEYINPUT90), .B1(new_n216), .B2(new_n679), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(KEYINPUT90), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  OR2_X1    g0484(.A1(new_n643), .A2(new_n644), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n653), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n651), .B1(new_n642), .B2(new_n650), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n663), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT29), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n655), .A2(new_n663), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(KEYINPUT29), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n639), .A2(new_n589), .A3(new_n299), .A4(new_n303), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT92), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n309), .A2(new_n695), .A3(new_n589), .A4(new_n639), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n518), .A2(new_n519), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n587), .B1(new_n698), .B2(new_n292), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n698), .A2(new_n313), .A3(new_n587), .A4(new_n617), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n697), .A2(new_n619), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT91), .A3(new_n313), .A4(new_n587), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n700), .A2(KEYINPUT93), .A3(new_n707), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n701), .A2(new_n704), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n664), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n700), .A2(new_n707), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n663), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n563), .A2(new_n324), .A3(new_n627), .A4(new_n664), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(KEYINPUT94), .A3(new_n714), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n716), .A2(new_n721), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n692), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n684), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(new_n261), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n206), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n678), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n669), .B2(G330), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n669), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n213), .B1(G20), .B2(new_n250), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n677), .A2(new_n348), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G45), .B2(new_n216), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n248), .B2(G45), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n677), .A2(new_n463), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G355), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G116), .B2(new_n210), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n738), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(new_n731), .ZN(new_n746));
  INV_X1    g0546(.A(new_n737), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n589), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G190), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G58), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(G190), .A3(new_n415), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n348), .B1(new_n750), .B2(new_n350), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n207), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n598), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n358), .A3(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n422), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n748), .A2(new_n358), .A3(G200), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n358), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n207), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n759), .B1(new_n372), .B2(new_n760), .C1(new_n252), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n753), .B(new_n763), .C1(G50), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n754), .A2(new_n749), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT96), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT96), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n457), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n769), .A2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n463), .B1(new_n750), .B2(new_n779), .C1(new_n780), .C2(new_n752), .ZN(new_n781));
  INV_X1    g0581(.A(new_n762), .ZN(new_n782));
  INV_X1    g0582(.A(new_n755), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(G294), .B1(new_n783), .B2(G303), .ZN(new_n784));
  INV_X1    g0584(.A(new_n760), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n784), .B(new_n789), .C1(new_n790), .C2(new_n757), .ZN(new_n791));
  INV_X1    g0591(.A(new_n774), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n781), .B(new_n791), .C1(G329), .C2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n770), .A2(new_n777), .B1(new_n778), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n736), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n746), .B1(new_n747), .B2(new_n794), .C1(new_n669), .C2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n733), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  NOR2_X1   g0598(.A1(new_n437), .A2(new_n663), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n438), .A2(new_n439), .B1(new_n435), .B2(new_n664), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n437), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n691), .B(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n731), .B1(new_n805), .B2(new_n725), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n725), .B2(new_n805), .ZN(new_n807));
  INV_X1    g0607(.A(new_n731), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n747), .A2(new_n735), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT98), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n808), .B1(new_n811), .B2(new_n350), .ZN(new_n812));
  INV_X1    g0612(.A(new_n752), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n348), .B1(new_n813), .B2(G294), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n814), .B1(new_n256), .B2(new_n750), .C1(new_n774), .C2(new_n779), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n757), .A2(new_n598), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G97), .B2(new_n782), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n422), .B2(new_n755), .C1(new_n790), .C2(new_n760), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n818), .C1(G303), .C2(new_n769), .ZN(new_n819));
  INV_X1    g0619(.A(new_n750), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n813), .A2(G143), .B1(new_n820), .B2(G159), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n326), .B2(new_n760), .C1(new_n768), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n782), .A2(G58), .B1(new_n783), .B2(G50), .ZN(new_n826));
  INV_X1    g0626(.A(new_n757), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n463), .B1(new_n827), .B2(G68), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(new_n774), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n823), .B2(new_n824), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n819), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n812), .B1(new_n747), .B2(new_n832), .C1(new_n804), .C2(new_n735), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n807), .A2(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n728), .A2(new_n206), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n503), .B2(new_n661), .ZN(new_n837));
  INV_X1    g0637(.A(new_n661), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n484), .A2(KEYINPUT100), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n481), .B1(new_n503), .B2(new_n504), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n470), .B2(new_n499), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n443), .B1(new_n494), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n487), .B2(new_n838), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n481), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n846), .A2(new_n838), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n511), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT101), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n481), .B(KEYINPUT17), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n505), .A2(new_n488), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n840), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n840), .A2(new_n843), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n859), .B2(new_n844), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n854), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(new_n840), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n632), .B2(new_n483), .ZN(new_n863));
  INV_X1    g0663(.A(new_n844), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n841), .B1(new_n840), .B2(new_n843), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n853), .A2(KEYINPUT38), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n718), .A2(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n722), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n382), .A2(new_n664), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n413), .A2(new_n418), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n407), .A2(G169), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT14), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n410), .A3(new_n409), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n383), .B(new_n663), .C1(new_n877), .C2(new_n417), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n803), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT40), .B1(new_n869), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n852), .A2(new_n867), .ZN(new_n882));
  OAI211_X1 g0682(.A(KEYINPUT38), .B(new_n850), .C1(new_n511), .C2(new_n851), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  INV_X1    g0685(.A(new_n880), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n513), .A3(new_n871), .ZN(new_n889));
  AOI211_X1 g0689(.A(KEYINPUT40), .B(new_n880), .C1(new_n882), .C2(new_n883), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n860), .A2(new_n854), .A3(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT101), .B1(new_n866), .B2(new_n867), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n883), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n893), .B2(new_n886), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n513), .A2(new_n871), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(G330), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT102), .Z(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n804), .B(new_n664), .C1(new_n645), .C2(new_n654), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n800), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n874), .A2(new_n878), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT99), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n907), .A2(new_n884), .B1(new_n632), .B2(new_n661), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n877), .A2(new_n383), .A3(new_n664), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n634), .B1(new_n692), .B2(new_n512), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n835), .B1(new_n900), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n900), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n569), .A2(new_n567), .ZN(new_n920));
  INV_X1    g0720(.A(new_n568), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n922), .A2(KEYINPUT35), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(KEYINPUT35), .ZN(new_n924));
  NOR4_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(new_n256), .A4(new_n215), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT36), .Z(new_n926));
  OR3_X1    g0726(.A1(new_n216), .A2(new_n455), .A3(new_n350), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n201), .A2(G68), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(G1), .A3(new_n261), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n919), .A2(new_n926), .A3(new_n930), .ZN(G367));
  OAI211_X1 g0731(.A(new_n591), .B(new_n593), .C1(new_n577), .C2(new_n664), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n650), .A2(new_n663), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n563), .A2(new_n934), .A3(new_n671), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n591), .B1(new_n932), .B2(new_n560), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n664), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n605), .A2(new_n623), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n663), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n653), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT103), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n642), .A2(new_n940), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT104), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT104), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n938), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  MUX2_X1   g0749(.A(new_n948), .B(KEYINPUT43), .S(new_n946), .Z(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n938), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n934), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n670), .B2(new_n952), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n951), .A2(new_n670), .A3(new_n952), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n678), .B(KEYINPUT41), .Z(new_n955));
  INV_X1    g0755(.A(new_n670), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n675), .A2(new_n957), .A3(new_n934), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT45), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT106), .B1(new_n674), .B2(new_n952), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n674), .A2(new_n952), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n674), .A2(KEYINPUT44), .A3(new_n952), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n966), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(KEYINPUT107), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n956), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n958), .A2(new_n960), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT45), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n970), .A2(KEYINPUT107), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n968), .B2(new_n967), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n978), .A3(new_n670), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n672), .B1(new_n666), .B2(new_n671), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n669), .A2(KEYINPUT108), .A3(G330), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT108), .B1(new_n669), .B2(G330), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n980), .A2(new_n983), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n726), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT109), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT109), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n726), .A2(new_n984), .A3(new_n988), .A4(new_n985), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n972), .A2(new_n979), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n955), .B1(new_n990), .B2(new_n726), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n953), .B(new_n954), .C1(new_n991), .C2(new_n730), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n738), .B1(new_n210), .B2(new_n604), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n739), .B2(new_n234), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n769), .A2(G143), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n762), .A2(new_n372), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n760), .A2(new_n457), .B1(new_n757), .B2(new_n350), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G58), .C2(new_n783), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n792), .A2(G137), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n348), .B1(new_n752), .B2(new_n326), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n201), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n820), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n995), .A2(new_n998), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n827), .A2(G97), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n463), .B(new_n1004), .C1(new_n774), .C2(new_n786), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n769), .A2(G311), .ZN(new_n1007));
  INV_X1    g0807(.A(G294), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n760), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(G303), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n752), .A2(new_n1010), .B1(new_n750), .B2(new_n790), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G107), .C2(new_n782), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n755), .A2(new_n1013), .A3(new_n256), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n755), .B2(new_n256), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1007), .A2(new_n1012), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1003), .B1(new_n1006), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n808), .B(new_n994), .C1(new_n1020), .C2(new_n737), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n946), .B2(new_n795), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n992), .A2(new_n1022), .ZN(G387));
  AND2_X1   g0823(.A1(new_n984), .A2(new_n985), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n679), .B1(new_n1024), .B2(new_n726), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n726), .B2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n730), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n680), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n742), .A2(new_n1028), .B1(new_n422), .B2(new_n677), .ZN(new_n1029));
  INV_X1    g0829(.A(G45), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n239), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n331), .A2(G50), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT50), .Z(new_n1033));
  OAI211_X1 g0833(.A(new_n680), .B(new_n1030), .C1(new_n372), .C2(new_n350), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n739), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n808), .B1(new_n1036), .B2(new_n738), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n463), .B1(new_n820), .B2(G68), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n335), .B2(new_n752), .C1(new_n774), .C2(new_n326), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n782), .A2(new_n429), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(new_n1004), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n350), .B2(new_n755), .C1(new_n331), .C2(new_n760), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(G159), .C2(new_n769), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n813), .A2(G317), .B1(new_n820), .B2(G303), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n779), .B2(new_n760), .C1(new_n768), .C2(new_n780), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n782), .A2(G283), .B1(new_n783), .B2(G294), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1052));
  INV_X1    g0852(.A(G326), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n463), .B1(new_n256), .B2(new_n757), .C1(new_n774), .C2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1051), .B2(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1043), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1037), .B1(new_n747), .B2(new_n1056), .C1(new_n666), .C2(new_n795), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1027), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1026), .A2(new_n1058), .ZN(G393));
  INV_X1    g0859(.A(new_n979), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n670), .B1(new_n976), .B2(new_n978), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n986), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n678), .A3(new_n990), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n244), .A2(new_n677), .A3(new_n348), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n738), .B1(new_n252), .B2(new_n210), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n731), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n934), .A2(new_n795), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n768), .A2(new_n786), .B1(new_n779), .B2(new_n752), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  AOI211_X1 g0869(.A(new_n348), .B(new_n758), .C1(G294), .C2(new_n820), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n760), .A2(new_n1010), .B1(new_n755), .B2(new_n790), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G116), .B2(new_n782), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n780), .C2(new_n774), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n768), .A2(new_n326), .B1(new_n457), .B2(new_n752), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n348), .B1(new_n750), .B2(new_n331), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n816), .B(new_n1078), .C1(new_n792), .C2(G143), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n760), .A2(new_n201), .B1(new_n755), .B2(new_n372), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G77), .B2(new_n782), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1069), .A2(new_n1073), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT114), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1066), .B(new_n1067), .C1(new_n737), .C2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n730), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1087), .ZN(G390));
  AOI21_X1  g0888(.A(new_n912), .B1(new_n902), .B2(new_n903), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n910), .B2(new_n913), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n724), .A2(G330), .A3(new_n903), .A4(new_n804), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n799), .B1(new_n689), .B2(new_n802), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n903), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n911), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n869), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT115), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1089), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n861), .A2(new_n868), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n883), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1097), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n689), .A2(new_n802), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n800), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n912), .B1(new_n1104), .B2(new_n903), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n724), .A2(G330), .A3(new_n804), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1105), .A2(new_n893), .B1(new_n1107), .B2(new_n903), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1101), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n869), .A2(new_n1094), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1101), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n871), .A2(new_n879), .A3(G330), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1096), .A2(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n871), .A2(G330), .A3(new_n804), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1093), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1091), .A2(new_n1116), .A3(new_n1092), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1113), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n902), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND4_X1   g0920(.A1(G330), .A2(new_n441), .A3(new_n511), .A4(new_n871), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n916), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT116), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT116), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1114), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1120), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1114), .B2(KEYINPUT117), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1113), .B1(new_n1090), .B2(new_n1110), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1090), .A2(new_n1095), .A3(KEYINPUT115), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1102), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n678), .B(new_n1128), .C1(new_n1132), .C2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n735), .B1(new_n910), .B2(new_n913), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n348), .B1(new_n820), .B2(G97), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n256), .B2(new_n752), .C1(new_n774), .C2(new_n1008), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n756), .B1(G68), .B2(new_n827), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n350), .B2(new_n762), .C1(new_n422), .C2(new_n760), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G283), .C2(new_n769), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n782), .A2(G159), .B1(new_n827), .B2(new_n1001), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1146), .B1(new_n822), .B2(new_n760), .C1(new_n768), .C2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  AOI21_X1  g0949(.A(new_n463), .B1(new_n820), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1150), .B1(new_n829), .B2(new_n752), .C1(new_n774), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n783), .A2(G150), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT53), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1148), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n737), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n808), .B1(new_n811), .B2(new_n331), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1136), .A2(new_n729), .B1(new_n1140), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1139), .A2(new_n1160), .ZN(G378));
  NAND2_X1  g0961(.A1(new_n1128), .A2(new_n1122), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n338), .A2(new_n838), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n371), .B(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n888), .B2(G330), .ZN(new_n1168));
  OAI211_X1 g0968(.A(G330), .B(new_n1167), .C1(new_n890), .C2(new_n894), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n915), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1167), .ZN(new_n1172));
  INV_X1    g0972(.A(G330), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n895), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n908), .A2(new_n914), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n1169), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1163), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n679), .B1(new_n1162), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1168), .A2(new_n1170), .A3(new_n915), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1175), .B1(new_n1174), .B2(new_n1169), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1122), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1114), .B2(new_n1127), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1163), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n731), .B1(new_n1001), .B2(new_n809), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n348), .A2(G41), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n335), .B1(G33), .B2(G41), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1187), .B1(new_n752), .B2(new_n422), .C1(new_n604), .C2(new_n750), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n792), .B2(G283), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n760), .A2(new_n252), .B1(new_n757), .B2(new_n751), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n996), .B(new_n1192), .C1(G77), .C2(new_n783), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n256), .C2(new_n768), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1189), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n752), .A2(new_n1147), .B1(new_n750), .B2(new_n822), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G132), .B2(new_n785), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n782), .A2(G150), .B1(new_n783), .B2(new_n1149), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1151), .C2(new_n768), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n792), .A2(G124), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n827), .C2(G159), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1201), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1186), .B1(new_n1206), .B2(new_n737), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1167), .B2(new_n735), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT118), .Z(new_n1209));
  NAND2_X1  g1009(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n730), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1185), .A2(new_n1211), .ZN(G375));
  NAND2_X1  g1012(.A1(new_n1120), .A2(new_n730), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n731), .B1(new_n810), .B2(G68), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1040), .B1(new_n350), .B2(new_n757), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n774), .A2(new_n1010), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n760), .A2(new_n256), .B1(new_n755), .B2(new_n252), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n463), .B1(new_n750), .B2(new_n422), .C1(new_n790), .C2(new_n752), .ZN(new_n1218));
  OR4_X1    g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n768), .A2(new_n1008), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n768), .A2(new_n829), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n792), .A2(G128), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n782), .A2(G50), .B1(new_n827), .B2(G58), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n785), .A2(new_n1149), .B1(new_n783), .B2(G159), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n348), .B1(new_n752), .B2(new_n822), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n820), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1219), .A2(new_n1220), .B1(new_n1221), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1214), .B1(new_n1228), .B2(new_n737), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n903), .B2(new_n735), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1213), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1124), .A2(new_n1126), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n955), .ZN(G381));
  OAI21_X1  g1035(.A(new_n678), .B1(new_n1136), .B2(new_n1131), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT119), .B1(new_n1239), .B2(new_n1159), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT119), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1139), .A2(new_n1241), .A3(new_n1160), .ZN(new_n1242));
  AND4_X1   g1042(.A1(new_n1211), .A2(new_n1240), .A3(new_n1185), .A4(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1026), .A2(new_n797), .A3(new_n1058), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(G384), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(G407));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n662), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(new_n1248), .A3(G213), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT120), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n992), .A2(new_n1022), .A3(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT122), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT122), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n992), .A2(new_n1254), .A3(new_n1022), .A4(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(G390), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1244), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1252), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n992), .A2(KEYINPUT123), .A3(new_n1022), .A4(G390), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n1257), .A3(new_n1260), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1162), .A2(new_n1210), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1211), .B1(new_n1269), .B2(new_n955), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1240), .A2(new_n1242), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1185), .A2(G378), .A3(new_n1211), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT60), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n678), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1234), .B2(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1277), .B1(new_n1281), .B2(new_n1231), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1281), .A2(new_n1277), .A3(new_n1231), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AND4_X1   g1085(.A1(new_n1268), .A2(new_n1273), .A3(new_n1276), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1275), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1281), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G384), .A3(new_n1232), .ZN(new_n1290));
  INV_X1    g1090(.A(G2897), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1276), .A2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1290), .A2(new_n1282), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1290), .B2(new_n1282), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1287), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1286), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1285), .ZN(new_n1298));
  XOR2_X1   g1098(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1267), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT121), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n1283), .A2(new_n1284), .B1(new_n1291), .B2(new_n1276), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1290), .A2(new_n1282), .A3(new_n1292), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(KEYINPUT121), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1267), .B(new_n1287), .C1(new_n1307), .C2(new_n1288), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT63), .B1(new_n1288), .B2(new_n1285), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1308), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1251), .B1(new_n1301), .B2(new_n1312), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1288), .A2(new_n1295), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1288), .A2(new_n1268), .A3(new_n1285), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1300), .A2(new_n1314), .A3(new_n1287), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1267), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1309), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1320), .A3(KEYINPUT125), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1321), .ZN(G405));
  NOR2_X1   g1122(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(new_n1267), .B(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(G375), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1272), .A3(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1324), .B(new_n1327), .ZN(G402));
endmodule


