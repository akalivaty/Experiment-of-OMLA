//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT67), .A2(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT67), .A2(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G116), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT68), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(G119), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT2), .A2(G113), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT2), .A2(G113), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(new_n196), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT69), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n191), .A2(new_n196), .A3(new_n202), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n191), .A2(new_n196), .ZN(new_n205));
  INV_X1    g019(.A(new_n199), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT11), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n212), .B2(G134), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT64), .A3(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(KEYINPUT65), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT0), .A3(G128), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n229), .A3(G131), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n223), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n212), .A2(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n209), .A2(G137), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n221), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  INV_X1    g051(.A(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G143), .ZN(new_n239));
  INV_X1    g053(.A(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n236), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(new_n224), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n235), .A2(new_n244), .A3(new_n222), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT30), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n208), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n223), .A2(new_n228), .A3(new_n230), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT30), .B1(new_n249), .B2(new_n246), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n188), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n246), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n201), .A2(new_n203), .B1(new_n206), .B2(new_n205), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n246), .A2(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(new_n249), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n257), .A3(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n255), .A3(new_n246), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(KEYINPUT26), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(G101), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n261), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n260), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n251), .B2(new_n258), .ZN(new_n271));
  INV_X1    g085(.A(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT72), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n255), .B1(new_n249), .B2(new_n246), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT28), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n277), .A3(new_n272), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n252), .A2(new_n208), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n276), .B1(new_n284), .B2(new_n260), .ZN(new_n285));
  INV_X1    g099(.A(new_n277), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(KEYINPUT29), .A3(new_n272), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n187), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n268), .A2(new_n270), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n248), .A2(new_n188), .A3(new_n250), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT70), .B1(new_n254), .B2(new_n257), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT31), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n268), .B1(new_n285), .B2(new_n286), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n259), .A2(new_n299), .A3(new_n293), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n302), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT74), .B(G217), .Z(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G234), .B2(new_n290), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n189), .A2(new_n190), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n236), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT76), .B(G110), .ZN(new_n319));
  NOR2_X1   g133(.A1(G119), .A2(G128), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n315), .B2(G128), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n318), .B(new_n319), .C1(new_n322), .C2(new_n317), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT24), .B(G110), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(KEYINPUT77), .A3(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n333), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(G146), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT78), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n238), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n335), .A2(new_n341), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n332), .A2(new_n334), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n238), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n321), .A2(new_n324), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n318), .B1(new_n322), .B2(new_n317), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(G110), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT22), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(G137), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n340), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n338), .B1(new_n328), .B2(new_n329), .ZN(new_n358));
  INV_X1    g172(.A(new_n351), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n290), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n314), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n356), .A2(new_n360), .A3(new_n290), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n313), .A2(G902), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n360), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n311), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n304), .B2(new_n310), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT80), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n380), .A2(new_n383), .A3(new_n387), .A4(new_n384), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n390), .A3(G101), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n208), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n391), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT84), .B1(new_n255), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G113), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n189), .A2(G116), .A3(new_n190), .ZN(new_n398));
  XOR2_X1   g212(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n205), .B2(new_n399), .ZN(new_n401));
  INV_X1    g215(.A(new_n384), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n379), .A2(G107), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n388), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n204), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n394), .A2(new_n396), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G110), .B(G122), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT86), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n408), .B2(new_n410), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n396), .A2(new_n407), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n409), .A4(new_n394), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n394), .A2(new_n396), .A3(new_n409), .A4(new_n407), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT87), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(KEYINPUT6), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n352), .A2(G224), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT88), .Z(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT89), .Z(new_n425));
  OR2_X1    g239(.A1(new_n244), .A2(G125), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n227), .A2(G125), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n425), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n204), .A2(new_n401), .A3(new_n405), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n409), .B(KEYINPUT8), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n191), .A2(new_n196), .A3(KEYINPUT5), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n201), .A2(new_n203), .B1(new_n400), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n433), .C1(new_n405), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n426), .A2(new_n427), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n426), .B2(new_n427), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT90), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n418), .A2(new_n420), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n378), .B1(new_n431), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n415), .B2(new_n421), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n419), .B(new_n417), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n290), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  INV_X1    g267(.A(new_n378), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n377), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G113), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(new_n379), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n263), .A2(G214), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n240), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G131), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(G143), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n221), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(KEYINPUT17), .A3(G131), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(new_n347), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n331), .A2(new_n238), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n462), .A2(new_n469), .B1(new_n470), .B2(new_n337), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(KEYINPUT18), .A3(G131), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n458), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n458), .B(new_n473), .C1(new_n467), .C2(new_n347), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n290), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G475), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n331), .B(KEYINPUT19), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n461), .A2(new_n463), .B1(new_n480), .B2(new_n238), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(new_n336), .B1(new_n472), .B2(new_n471), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n475), .B1(new_n458), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n484), .A4(new_n485), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n479), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(G952), .A3(new_n352), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(G902), .A3(G953), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G128), .B(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT13), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n236), .A2(KEYINPUT13), .A3(G143), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n209), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n503), .B1(new_n209), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT92), .B1(new_n192), .B2(G122), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  INV_X1    g320(.A(G122), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(G116), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n193), .A2(new_n195), .A3(G122), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n509), .A2(new_n510), .A3(new_n382), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n382), .B1(new_n509), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT93), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n504), .B(new_n515), .C1(new_n512), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n500), .A2(new_n209), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n500), .A2(new_n209), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n510), .A2(KEYINPUT14), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n509), .B1(new_n510), .B2(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g336(.A(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT9), .B(G234), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n312), .A2(G953), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n514), .A2(new_n516), .B1(new_n523), .B2(new_n520), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT94), .B1(new_n531), .B2(new_n528), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n530), .B(new_n532), .C1(new_n525), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n290), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n536), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n533), .B2(new_n290), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n491), .A2(new_n499), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n456), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G469), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G140), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT81), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n352), .A2(G227), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n545), .B(new_n546), .Z(new_n547));
  AND2_X1   g361(.A1(new_n244), .A2(KEYINPUT10), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n392), .A2(new_n228), .B1(new_n406), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT82), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n236), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n239), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n224), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n242), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n406), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(KEYINPUT83), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT83), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n549), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n223), .A2(new_n230), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n549), .B(new_n562), .C1(new_n559), .C2(new_n560), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n547), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n556), .B1(new_n244), .B2(new_n406), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n563), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT12), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n565), .A2(new_n569), .A3(new_n547), .A4(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n543), .B(new_n290), .C1(new_n566), .C2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n543), .A2(new_n290), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n565), .A2(new_n571), .A3(new_n569), .ZN(new_n576));
  INV_X1    g390(.A(new_n547), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n564), .A2(new_n565), .A3(new_n547), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n573), .B(new_n575), .C1(new_n580), .C2(new_n543), .ZN(new_n581));
  OAI21_X1  g395(.A(G221), .B1(new_n527), .B2(G902), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n542), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n374), .A2(new_n376), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT95), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n387), .ZN(G3));
  NAND2_X1  g401(.A1(new_n534), .A2(new_n535), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT98), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n534), .A2(new_n590), .A3(new_n535), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n533), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n525), .A2(KEYINPUT96), .A3(new_n529), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n531), .B1(new_n595), .B2(new_n528), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(KEYINPUT33), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n594), .A2(new_n596), .A3(new_n599), .A4(KEYINPUT33), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n535), .A2(G902), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n593), .A2(new_n598), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n589), .A2(new_n591), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n489), .A2(new_n490), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n478), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n607));
  INV_X1    g421(.A(new_n377), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n431), .A2(new_n378), .A3(new_n449), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n454), .B1(new_n451), .B2(new_n453), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n606), .A2(new_n607), .A3(new_n611), .A4(new_n499), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n603), .A2(new_n499), .A3(new_n605), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT99), .B1(new_n613), .B2(new_n456), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT71), .B1(new_n301), .B2(new_n302), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n301), .A2(new_n290), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n619), .A2(new_n187), .ZN(new_n620));
  AND4_X1   g434(.A1(new_n618), .A2(new_n620), .A3(new_n371), .A4(new_n583), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n540), .ZN(new_n625));
  INV_X1    g439(.A(new_n486), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n487), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n479), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n611), .A2(new_n499), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NAND2_X1  g447(.A1(new_n620), .A2(new_n618), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n340), .A2(new_n351), .A3(new_n635), .ZN(new_n636));
  OAI22_X1  g450(.A1(new_n358), .A2(new_n359), .B1(KEYINPUT36), .B2(new_n357), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n368), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n367), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n581), .A3(new_n582), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n542), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT37), .B(G110), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(new_n641), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT32), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n301), .A2(KEYINPUT32), .A3(new_n302), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n289), .A2(new_n290), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n272), .B1(new_n259), .B2(new_n260), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n280), .B1(new_n651), .B2(new_n262), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n650), .B1(new_n652), .B2(new_n273), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n649), .B1(new_n653), .B2(new_n187), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n611), .B(new_n647), .C1(new_n648), .C2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT101), .B(G900), .Z(new_n656));
  AOI21_X1  g470(.A(new_n494), .B1(new_n656), .B2(new_n496), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n478), .B(new_n658), .C1(new_n626), .C2(new_n487), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n540), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n655), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n641), .B1(new_n304), .B2(new_n310), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n663), .A2(new_n660), .A3(new_n664), .A4(new_n611), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n261), .A2(new_n272), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n270), .A2(new_n274), .ZN(new_n669));
  AOI21_X1  g483(.A(G902), .B1(new_n669), .B2(new_n268), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n187), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n303), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n310), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT103), .Z(new_n674));
  XOR2_X1   g488(.A(new_n657), .B(KEYINPUT39), .Z(new_n675));
  NAND2_X1  g489(.A1(new_n583), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n609), .A2(new_n610), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n640), .A2(new_n491), .A3(new_n608), .A4(new_n540), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n674), .A2(new_n677), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT104), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n603), .A2(new_n605), .A3(new_n658), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n603), .A2(new_n686), .A3(new_n605), .A4(new_n658), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n655), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n238), .ZN(G48));
  OAI21_X1  g504(.A(new_n290), .B1(new_n566), .B2(new_n572), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n573), .ZN(new_n693));
  INV_X1    g507(.A(new_n582), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n615), .A2(new_n375), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n371), .B(new_n695), .C1(new_n648), .C2(new_n654), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n699), .B1(new_n700), .B2(new_n629), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n375), .A2(new_n630), .A3(KEYINPUT106), .A4(new_n695), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NAND2_X1  g518(.A1(new_n695), .A2(new_n611), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n638), .B1(new_n363), .B2(new_n366), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n541), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n311), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND4_X1  g524(.A1(new_n678), .A2(new_n377), .A3(new_n625), .A4(new_n605), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n611), .A2(KEYINPUT107), .A3(new_n625), .A4(new_n605), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n619), .A2(new_n187), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n692), .A2(new_n499), .A3(new_n582), .A4(new_n573), .ZN(new_n717));
  INV_X1    g531(.A(new_n302), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n297), .A2(new_n300), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n287), .A2(new_n288), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n268), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n716), .A2(new_n370), .A3(new_n717), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n715), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR2_X1   g539(.A1(new_n722), .A2(new_n707), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n620), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n688), .A2(new_n705), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n333), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n579), .B1(new_n578), .B2(KEYINPUT108), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n576), .B2(new_n577), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n733), .A3(new_n543), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n573), .A2(new_n575), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n582), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n609), .A2(new_n610), .A3(new_n377), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n375), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n730), .B1(new_n739), .B2(new_n688), .ZN(new_n740));
  INV_X1    g554(.A(new_n688), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n305), .A2(new_n308), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n370), .B1(new_n304), .B2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(KEYINPUT42), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NOR2_X1   g560(.A1(new_n739), .A2(new_n661), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n209), .ZN(G36));
  NAND2_X1  g562(.A1(new_n603), .A2(new_n491), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT43), .Z(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n634), .A3(new_n640), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT109), .Z(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n731), .A2(new_n755), .A3(new_n733), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n543), .B1(new_n580), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n574), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n573), .B1(new_n758), .B2(KEYINPUT46), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n582), .B(new_n675), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n737), .B1(new_n751), .B2(new_n752), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  OAI21_X1  g579(.A(new_n582), .B1(new_n759), .B2(new_n760), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT47), .Z(new_n767));
  NOR3_X1   g581(.A1(new_n311), .A2(new_n371), .A3(new_n737), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n741), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(new_n674), .ZN(new_n771));
  INV_X1    g585(.A(new_n679), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n693), .B(KEYINPUT49), .Z(new_n773));
  NOR4_X1   g587(.A1(new_n749), .A2(new_n370), .A3(new_n608), .A4(new_n694), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n701), .A2(new_n702), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n696), .A2(new_n709), .A3(new_n724), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT110), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n700), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n311), .A2(new_n708), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n780), .A2(new_n615), .B1(new_n781), .B2(new_n706), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n703), .A3(new_n783), .A4(new_n724), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n540), .A2(new_n628), .A3(new_n658), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n737), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT111), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n785), .B2(new_n737), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n311), .A3(new_n647), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n716), .A2(new_n707), .A3(new_n722), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n687), .A3(new_n685), .A4(new_n738), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n603), .A2(new_n491), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n491), .A2(new_n540), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n611), .A2(new_n795), .A3(new_n499), .A4(new_n796), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n621), .A2(new_n797), .B1(new_n642), .B2(new_n542), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n585), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n747), .B1(new_n740), .B2(new_n744), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n779), .A2(new_n784), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n728), .B1(new_n662), .B2(new_n665), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n641), .B(new_n456), .C1(new_n304), .C2(new_n310), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n638), .B(new_n657), .C1(new_n363), .C2(new_n366), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(new_n582), .C1(new_n735), .C2(new_n734), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n310), .B2(new_n672), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n803), .A2(new_n741), .B1(new_n715), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n802), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n776), .B1(new_n801), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n728), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n666), .A2(new_n812), .A3(new_n807), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n777), .A2(new_n778), .ZN(new_n818));
  INV_X1    g632(.A(new_n747), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n745), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n585), .A2(new_n794), .A3(new_n798), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT54), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n817), .A2(new_n779), .A3(new_n784), .A4(new_n822), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n776), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(KEYINPUT54), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n750), .A2(new_n494), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n829), .A2(new_n370), .A3(new_n716), .A4(new_n722), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n608), .A3(new_n772), .A4(new_n695), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT50), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n831), .B(new_n833), .Z(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n832), .B2(KEYINPUT50), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n693), .A2(new_n582), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n787), .B(new_n830), .C1(new_n767), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n787), .A2(new_n695), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT113), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n370), .A2(new_n493), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n771), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n605), .A3(new_n603), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n839), .A2(new_n494), .A3(new_n750), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n792), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n743), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n850), .A2(KEYINPUT48), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n352), .A2(G952), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n830), .B2(new_n706), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n849), .B2(new_n851), .ZN(new_n856));
  INV_X1    g670(.A(new_n841), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n853), .B(new_n856), .C1(new_n606), .C2(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n828), .A2(new_n847), .A3(new_n848), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(G952), .A2(G953), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n775), .B1(new_n859), .B2(new_n860), .ZN(G75));
  NOR2_X1   g675(.A1(new_n352), .A2(G952), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AND4_X1   g677(.A1(KEYINPUT53), .A2(new_n818), .A3(new_n799), .A4(new_n800), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n826), .A2(new_n776), .B1(new_n817), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n290), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT56), .B1(new_n866), .B2(G210), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n422), .A2(new_n430), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n451), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT115), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT55), .Z(new_n871));
  OAI21_X1  g685(.A(new_n863), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n867), .B2(new_n871), .ZN(G51));
  XNOR2_X1  g687(.A(new_n865), .B(KEYINPUT54), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n574), .B(KEYINPUT57), .Z(new_n875));
  OAI22_X1  g689(.A1(new_n874), .A2(new_n875), .B1(new_n566), .B2(new_n572), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n756), .A2(new_n757), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT116), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n866), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n862), .B1(new_n876), .B2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  INV_X1    g695(.A(new_n483), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n862), .ZN(G60));
  NAND3_X1  g699(.A1(new_n593), .A2(new_n600), .A3(new_n598), .ZN(new_n886));
  XNOR2_X1  g700(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n535), .A2(new_n290), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n863), .B1(new_n874), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n886), .B1(new_n828), .B2(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G63));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT60), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n865), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n356), .A2(new_n360), .ZN(new_n903));
  INV_X1    g717(.A(new_n901), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n824), .A2(KEYINPUT119), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n863), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n636), .A2(new_n637), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT119), .B1(new_n824), .B2(new_n904), .ZN(new_n909));
  AOI211_X1 g723(.A(new_n899), .B(new_n901), .C1(new_n811), .C2(new_n823), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n902), .A2(new_n905), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n908), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n907), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n898), .B1(new_n916), .B2(KEYINPUT61), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n909), .A2(new_n910), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n862), .B1(new_n918), .B2(new_n903), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n913), .B2(new_n908), .ZN(new_n920));
  INV_X1    g734(.A(new_n908), .ZN(new_n921));
  AOI211_X1 g735(.A(KEYINPUT120), .B(new_n921), .C1(new_n902), .C2(new_n905), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(KEYINPUT121), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n917), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n919), .B(KEYINPUT61), .C1(new_n920), .C2(new_n922), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n912), .A2(new_n915), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n919), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n932), .ZN(G66));
  NAND2_X1  g747(.A1(G224), .A2(G953), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n497), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n779), .A2(new_n784), .A3(new_n585), .A4(new_n798), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT123), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n352), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n415), .B(new_n421), .C1(G898), .C2(new_n352), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  OAI21_X1  g754(.A(new_n254), .B1(new_n231), .B2(new_n247), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(new_n480), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n795), .A2(new_n796), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n676), .A3(new_n737), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n374), .A2(new_n376), .A3(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n764), .A2(new_n769), .A3(new_n947), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n689), .B(new_n728), .C1(new_n665), .C2(new_n662), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n682), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n944), .B1(new_n956), .B2(new_n352), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n352), .B1(G227), .B2(G900), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n942), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n762), .A2(new_n715), .A3(new_n743), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n764), .A2(new_n769), .A3(new_n949), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n800), .B(KEYINPUT126), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n963), .B1(new_n969), .B2(new_n352), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n958), .A2(new_n960), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n959), .B1(new_n957), .B2(new_n970), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n969), .B2(new_n937), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n978), .A2(new_n272), .A3(new_n261), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n954), .A2(new_n937), .A3(new_n955), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n668), .B1(new_n980), .B2(new_n976), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n269), .A2(new_n296), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n982), .B2(new_n273), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n827), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n863), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n979), .A2(new_n981), .A3(new_n985), .ZN(G57));
endmodule


