

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(KEYINPUT102), .ZN(n670) );
  XNOR2_X1 U550 ( .A(n670), .B(KEYINPUT29), .ZN(n671) );
  XNOR2_X1 U551 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U552 ( .A1(G651), .A2(G543), .ZN(n787) );
  NOR2_X2 U553 ( .A1(G2105), .A2(n525), .ZN(n877) );
  NAND2_X1 U554 ( .A1(G85), .A2(n787), .ZN(n515) );
  XOR2_X1 U555 ( .A(KEYINPUT0), .B(G543), .Z(n576) );
  INV_X1 U556 ( .A(G651), .ZN(n516) );
  NOR2_X1 U557 ( .A1(n576), .A2(n516), .ZN(n788) );
  NAND2_X1 U558 ( .A1(G72), .A2(n788), .ZN(n514) );
  NAND2_X1 U559 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X1 U560 ( .A1(G543), .A2(n516), .ZN(n518) );
  XNOR2_X1 U561 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n517) );
  XNOR2_X1 U562 ( .A(n518), .B(n517), .ZN(n781) );
  NAND2_X1 U563 ( .A1(G60), .A2(n781), .ZN(n521) );
  NOR2_X1 U564 ( .A1(G651), .A2(n576), .ZN(n519) );
  XOR2_X1 U565 ( .A(KEYINPUT65), .B(n519), .Z(n783) );
  NAND2_X1 U566 ( .A1(G47), .A2(n783), .ZN(n520) );
  NAND2_X1 U567 ( .A1(n521), .A2(n520), .ZN(n522) );
  OR2_X1 U568 ( .A1(n523), .A2(n522), .ZN(G290) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n524), .Z(n876) );
  AND2_X1 U571 ( .A1(G138), .A2(n876), .ZN(n531) );
  INV_X1 U572 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G102), .A2(n877), .ZN(n529) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U575 ( .A1(G114), .A2(n872), .ZN(n527) );
  AND2_X1 U576 ( .A1(n525), .A2(G2105), .ZN(n873) );
  NAND2_X1 U577 ( .A1(G126), .A2(n873), .ZN(n526) );
  AND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U580 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U581 ( .A1(G125), .A2(n873), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n532), .B(KEYINPUT66), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G101), .A2(n877), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G137), .A2(n876), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G113), .A2(n872), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U589 ( .A1(n539), .A2(n538), .ZN(G160) );
  NAND2_X1 U590 ( .A1(G64), .A2(n781), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G52), .A2(n783), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U593 ( .A1(G90), .A2(n787), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G77), .A2(n788), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U597 ( .A1(n546), .A2(n545), .ZN(G171) );
  INV_X1 U598 ( .A(G171), .ZN(G301) );
  NAND2_X1 U599 ( .A1(G65), .A2(n781), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G53), .A2(n783), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT68), .B(n549), .Z(n553) );
  NAND2_X1 U603 ( .A1(G91), .A2(n787), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G78), .A2(n788), .ZN(n550) );
  AND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(G299) );
  XOR2_X1 U607 ( .A(KEYINPUT4), .B(KEYINPUT76), .Z(n555) );
  NAND2_X1 U608 ( .A1(G89), .A2(n787), .ZN(n554) );
  XNOR2_X1 U609 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U610 ( .A(KEYINPUT75), .B(n556), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n788), .A2(G76), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n559), .B(KEYINPUT5), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G63), .A2(n781), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G51), .A2(n783), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U618 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U619 ( .A(n565), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U620 ( .A1(G88), .A2(n787), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G75), .A2(n788), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n781), .A2(G62), .ZN(n568) );
  XOR2_X1 U624 ( .A(KEYINPUT84), .B(n568), .Z(n569) );
  NOR2_X1 U625 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n783), .A2(G50), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n572), .A2(n571), .ZN(G303) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G49), .A2(n783), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G74), .A2(G651), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U632 ( .A1(n781), .A2(n575), .ZN(n578) );
  NAND2_X1 U633 ( .A1(n576), .A2(G87), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U635 ( .A1(G73), .A2(n788), .ZN(n579) );
  XNOR2_X1 U636 ( .A(n579), .B(KEYINPUT2), .ZN(n586) );
  NAND2_X1 U637 ( .A1(G61), .A2(n781), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G48), .A2(n783), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G86), .A2(n787), .ZN(n582) );
  XNOR2_X1 U641 ( .A(KEYINPUT83), .B(n582), .ZN(n583) );
  NOR2_X1 U642 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(G305) );
  XNOR2_X1 U644 ( .A(G1986), .B(G290), .ZN(n969) );
  NOR2_X1 U645 ( .A1(G164), .A2(G1384), .ZN(n617) );
  NAND2_X1 U646 ( .A1(G160), .A2(G40), .ZN(n618) );
  NOR2_X1 U647 ( .A1(n617), .A2(n618), .ZN(n752) );
  NAND2_X1 U648 ( .A1(n969), .A2(n752), .ZN(n740) );
  NAND2_X1 U649 ( .A1(G131), .A2(n876), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G107), .A2(n872), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G95), .A2(n877), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT89), .B(n589), .ZN(n590) );
  NOR2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U655 ( .A1(n873), .A2(G119), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n863) );
  NAND2_X1 U657 ( .A1(G1991), .A2(n863), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT90), .B(n594), .Z(n603) );
  NAND2_X1 U659 ( .A1(G141), .A2(n876), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G117), .A2(n872), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n877), .A2(G105), .ZN(n597) );
  XOR2_X1 U663 ( .A(KEYINPUT38), .B(n597), .Z(n598) );
  NOR2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n873), .A2(G129), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n883) );
  AND2_X1 U667 ( .A1(G1996), .A2(n883), .ZN(n602) );
  NOR2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n927) );
  XNOR2_X1 U669 ( .A(KEYINPUT91), .B(n752), .ZN(n604) );
  NOR2_X1 U670 ( .A1(n927), .A2(n604), .ZN(n744) );
  XOR2_X1 U671 ( .A(KEYINPUT92), .B(n744), .Z(n616) );
  XNOR2_X1 U672 ( .A(G2067), .B(KEYINPUT37), .ZN(n605) );
  XOR2_X1 U673 ( .A(n605), .B(KEYINPUT87), .Z(n749) );
  NAND2_X1 U674 ( .A1(n873), .A2(G128), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n606), .B(KEYINPUT88), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G116), .A2(n872), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n609), .B(KEYINPUT35), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G140), .A2(n876), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G104), .A2(n877), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U682 ( .A(KEYINPUT34), .B(n612), .Z(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U684 ( .A(n615), .B(KEYINPUT36), .Z(n869) );
  NOR2_X1 U685 ( .A1(n749), .A2(n869), .ZN(n920) );
  NAND2_X1 U686 ( .A1(n752), .A2(n920), .ZN(n747) );
  NAND2_X1 U687 ( .A1(n616), .A2(n747), .ZN(n738) );
  XNOR2_X1 U688 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n694) );
  XOR2_X1 U689 ( .A(KEYINPUT25), .B(G2078), .Z(n943) );
  INV_X1 U690 ( .A(n617), .ZN(n619) );
  NOR2_X2 U691 ( .A1(n619), .A2(n618), .ZN(n656) );
  INV_X1 U692 ( .A(n656), .ZN(n684) );
  NOR2_X1 U693 ( .A1(n943), .A2(n684), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n620), .B(KEYINPUT96), .ZN(n622) );
  XOR2_X1 U695 ( .A(G1961), .B(KEYINPUT95), .Z(n1011) );
  NOR2_X1 U696 ( .A1(n656), .A2(n1011), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n675) );
  NOR2_X1 U698 ( .A1(n675), .A2(G301), .ZN(n623) );
  XOR2_X1 U699 ( .A(KEYINPUT97), .B(n623), .Z(n674) );
  NAND2_X1 U700 ( .A1(n787), .A2(G81), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT12), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G68), .A2(n788), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n627) );
  XNOR2_X1 U705 ( .A(n628), .B(n627), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n781), .A2(G56), .ZN(n629) );
  XOR2_X1 U707 ( .A(KEYINPUT14), .B(n629), .Z(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n783), .A2(G43), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n965) );
  NAND2_X1 U711 ( .A1(G1341), .A2(n684), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT99), .ZN(n638) );
  XOR2_X1 U713 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n636) );
  AND2_X1 U714 ( .A1(G1996), .A2(n656), .ZN(n635) );
  XOR2_X1 U715 ( .A(n636), .B(n635), .Z(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U717 ( .A(n639), .B(KEYINPUT100), .Z(n640) );
  NOR2_X1 U718 ( .A1(n965), .A2(n640), .ZN(n654) );
  NAND2_X1 U719 ( .A1(G1348), .A2(n684), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G2067), .A2(n656), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n660) );
  NAND2_X1 U722 ( .A1(n787), .A2(G92), .ZN(n643) );
  XOR2_X1 U723 ( .A(KEYINPUT71), .B(n643), .Z(n645) );
  NAND2_X1 U724 ( .A1(n781), .A2(G66), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U726 ( .A(KEYINPUT72), .B(n646), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G79), .A2(n788), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G54), .A2(n783), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U730 ( .A(KEYINPUT73), .B(n649), .Z(n650) );
  NOR2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U732 ( .A(KEYINPUT15), .B(n652), .Z(n984) );
  INV_X1 U733 ( .A(n984), .ZN(n889) );
  NAND2_X1 U734 ( .A1(n660), .A2(n889), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(n664) );
  NAND2_X1 U736 ( .A1(G1956), .A2(n684), .ZN(n655) );
  XNOR2_X1 U737 ( .A(KEYINPUT98), .B(n655), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n656), .A2(G2072), .ZN(n657) );
  XOR2_X1 U739 ( .A(KEYINPUT27), .B(n657), .Z(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n666) );
  NOR2_X1 U741 ( .A1(G299), .A2(n666), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n660), .A2(n889), .ZN(n661) );
  NOR2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U745 ( .A(KEYINPUT101), .B(n665), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G299), .A2(n666), .ZN(n667) );
  XOR2_X1 U747 ( .A(n667), .B(KEYINPUT28), .Z(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n696) );
  AND2_X1 U750 ( .A1(G301), .A2(n675), .ZN(n682) );
  NOR2_X1 U751 ( .A1(G2084), .A2(n684), .ZN(n699) );
  NAND2_X1 U752 ( .A1(G8), .A2(n684), .ZN(n733) );
  NOR2_X1 U753 ( .A1(G1966), .A2(n733), .ZN(n676) );
  XOR2_X1 U754 ( .A(KEYINPUT94), .B(n676), .Z(n697) );
  NAND2_X1 U755 ( .A1(G8), .A2(n697), .ZN(n677) );
  NOR2_X1 U756 ( .A1(n699), .A2(n677), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n678) );
  XNOR2_X1 U758 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U759 ( .A1(G168), .A2(n680), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U761 ( .A(n683), .B(KEYINPUT31), .ZN(n695) );
  NOR2_X1 U762 ( .A1(G1971), .A2(n733), .ZN(n686) );
  NOR2_X1 U763 ( .A1(G2090), .A2(n684), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n687) );
  AND2_X1 U765 ( .A1(G303), .A2(n687), .ZN(n689) );
  OR2_X1 U766 ( .A1(n695), .A2(n689), .ZN(n688) );
  OR2_X1 U767 ( .A1(n696), .A2(n688), .ZN(n691) );
  OR2_X1 U768 ( .A1(n689), .A2(G286), .ZN(n690) );
  AND2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U770 ( .A1(n692), .A2(G8), .ZN(n693) );
  XNOR2_X1 U771 ( .A(n694), .B(n693), .ZN(n721) );
  OR2_X1 U772 ( .A1(n696), .A2(n695), .ZN(n698) );
  AND2_X1 U773 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U774 ( .A1(n699), .A2(G8), .ZN(n700) );
  NAND2_X1 U775 ( .A1(n701), .A2(n700), .ZN(n715) );
  NOR2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U777 ( .A1(n974), .A2(KEYINPUT33), .ZN(n702) );
  NOR2_X1 U778 ( .A1(n702), .A2(n733), .ZN(n704) );
  XOR2_X1 U779 ( .A(G1981), .B(G305), .Z(n970) );
  INV_X1 U780 ( .A(n970), .ZN(n703) );
  NOR2_X1 U781 ( .A1(n704), .A2(n703), .ZN(n716) );
  AND2_X1 U782 ( .A1(n716), .A2(KEYINPUT33), .ZN(n708) );
  OR2_X1 U783 ( .A1(n708), .A2(n733), .ZN(n706) );
  AND2_X1 U784 ( .A1(n715), .A2(n706), .ZN(n705) );
  NAND2_X1 U785 ( .A1(n721), .A2(n705), .ZN(n714) );
  INV_X1 U786 ( .A(n706), .ZN(n712) );
  NOR2_X1 U787 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U788 ( .A1(G8), .A2(n707), .ZN(n710) );
  INV_X1 U789 ( .A(n708), .ZN(n709) );
  AND2_X1 U790 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U791 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n730) );
  NAND2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n975) );
  AND2_X1 U794 ( .A1(n715), .A2(n975), .ZN(n719) );
  INV_X1 U795 ( .A(n716), .ZN(n717) );
  OR2_X1 U796 ( .A1(n733), .A2(n717), .ZN(n726) );
  INV_X1 U797 ( .A(n726), .ZN(n718) );
  AND2_X1 U798 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n728) );
  INV_X1 U800 ( .A(n975), .ZN(n724) );
  NOR2_X1 U801 ( .A1(G1971), .A2(G303), .ZN(n722) );
  NOR2_X1 U802 ( .A1(n974), .A2(n722), .ZN(n723) );
  OR2_X1 U803 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U804 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U806 ( .A1(n730), .A2(n729), .ZN(n736) );
  NOR2_X1 U807 ( .A1(G1981), .A2(G305), .ZN(n731) );
  XNOR2_X1 U808 ( .A(n731), .B(KEYINPUT93), .ZN(n732) );
  XNOR2_X1 U809 ( .A(n732), .B(KEYINPUT24), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n755) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n883), .ZN(n917) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n863), .ZN(n924) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n741) );
  XOR2_X1 U817 ( .A(n741), .B(KEYINPUT105), .Z(n742) );
  NOR2_X1 U818 ( .A1(n924), .A2(n742), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n917), .A2(n745), .ZN(n746) );
  XNOR2_X1 U821 ( .A(KEYINPUT39), .B(n746), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n751) );
  AND2_X1 U823 ( .A1(n749), .A2(n869), .ZN(n750) );
  XOR2_X1 U824 ( .A(KEYINPUT106), .B(n750), .Z(n933) );
  NAND2_X1 U825 ( .A1(n751), .A2(n933), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U830 ( .A1(G135), .A2(n876), .ZN(n758) );
  NAND2_X1 U831 ( .A1(G111), .A2(n872), .ZN(n757) );
  NAND2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n761) );
  NAND2_X1 U833 ( .A1(n873), .A2(G123), .ZN(n759) );
  XOR2_X1 U834 ( .A(KEYINPUT18), .B(n759), .Z(n760) );
  NOR2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n877), .A2(G99), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n921) );
  XNOR2_X1 U838 ( .A(G2096), .B(n921), .ZN(n764) );
  OR2_X1 U839 ( .A1(G2100), .A2(n764), .ZN(G156) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  INV_X1 U841 ( .A(G82), .ZN(G220) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XOR2_X1 U843 ( .A(n765), .B(KEYINPUT10), .Z(n915) );
  NAND2_X1 U844 ( .A1(n915), .A2(G567), .ZN(n766) );
  XOR2_X1 U845 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U846 ( .A(G860), .ZN(n774) );
  OR2_X1 U847 ( .A1(n965), .A2(n774), .ZN(G153) );
  INV_X1 U848 ( .A(G868), .ZN(n806) );
  NOR2_X1 U849 ( .A1(G301), .A2(n806), .ZN(n768) );
  NOR2_X1 U850 ( .A1(G868), .A2(n889), .ZN(n767) );
  NOR2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U852 ( .A(KEYINPUT74), .B(n769), .ZN(G284) );
  NOR2_X1 U853 ( .A1(G286), .A2(n806), .ZN(n770) );
  XOR2_X1 U854 ( .A(KEYINPUT77), .B(n770), .Z(n773) );
  NOR2_X1 U855 ( .A1(G868), .A2(G299), .ZN(n771) );
  XNOR2_X1 U856 ( .A(KEYINPUT78), .B(n771), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n775), .A2(n984), .ZN(n776) );
  XNOR2_X1 U860 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n965), .ZN(n777) );
  XOR2_X1 U862 ( .A(KEYINPUT79), .B(n777), .Z(n780) );
  NAND2_X1 U863 ( .A1(G868), .A2(n984), .ZN(n778) );
  NOR2_X1 U864 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U866 ( .A1(n781), .A2(G67), .ZN(n782) );
  XOR2_X1 U867 ( .A(KEYINPUT81), .B(n782), .Z(n785) );
  NAND2_X1 U868 ( .A1(n783), .A2(G55), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U870 ( .A(KEYINPUT82), .B(n786), .ZN(n792) );
  NAND2_X1 U871 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U872 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n790), .A2(n789), .ZN(n791) );
  OR2_X1 U874 ( .A1(n792), .A2(n791), .ZN(n805) );
  NAND2_X1 U875 ( .A1(G559), .A2(n984), .ZN(n793) );
  XNOR2_X1 U876 ( .A(n793), .B(KEYINPUT80), .ZN(n803) );
  XNOR2_X1 U877 ( .A(n803), .B(n965), .ZN(n794) );
  NOR2_X1 U878 ( .A1(G860), .A2(n794), .ZN(n795) );
  XOR2_X1 U879 ( .A(n805), .B(n795), .Z(G145) );
  XOR2_X1 U880 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n796) );
  XNOR2_X1 U881 ( .A(G288), .B(n796), .ZN(n799) );
  XOR2_X1 U882 ( .A(G303), .B(G290), .Z(n797) );
  XNOR2_X1 U883 ( .A(n797), .B(n965), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n799), .B(n798), .ZN(n801) );
  XOR2_X1 U885 ( .A(G305), .B(n805), .Z(n800) );
  XNOR2_X1 U886 ( .A(n801), .B(n800), .ZN(n802) );
  XOR2_X1 U887 ( .A(n802), .B(G299), .Z(n890) );
  XNOR2_X1 U888 ( .A(n890), .B(n803), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n804), .A2(G868), .ZN(n808) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U897 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U898 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U899 ( .A1(G220), .A2(G219), .ZN(n813) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n813), .Z(n814) );
  XNOR2_X1 U901 ( .A(n814), .B(KEYINPUT86), .ZN(n815) );
  NOR2_X1 U902 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G96), .A2(n816), .ZN(n825) );
  NAND2_X1 U904 ( .A1(n825), .A2(G2106), .ZN(n820) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n817) );
  NOR2_X1 U906 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G108), .A2(n818), .ZN(n826) );
  NAND2_X1 U908 ( .A1(n826), .A2(G567), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n827) );
  NAND2_X1 U910 ( .A1(G661), .A2(G483), .ZN(n821) );
  NOR2_X1 U911 ( .A1(n827), .A2(n821), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n915), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  INV_X1 U923 ( .A(n827), .ZN(G319) );
  XNOR2_X1 U924 ( .A(G1986), .B(G2474), .ZN(n837) );
  XOR2_X1 U925 ( .A(G1981), .B(G1966), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1971), .B(G1961), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U928 ( .A(G1976), .B(G1956), .Z(n831) );
  XNOR2_X1 U929 ( .A(G1996), .B(G1991), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(G229) );
  XOR2_X1 U935 ( .A(KEYINPUT111), .B(G2084), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n840), .B(G2100), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2078), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(G227) );
  NAND2_X1 U945 ( .A1(G124), .A2(n873), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n872), .A2(G112), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U949 ( .A1(G136), .A2(n876), .ZN(n851) );
  NAND2_X1 U950 ( .A1(G100), .A2(n877), .ZN(n850) );
  NAND2_X1 U951 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U952 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U953 ( .A1(G139), .A2(n876), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G103), .A2(n877), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G115), .A2(n872), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G127), .A2(n873), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT47), .B(n858), .ZN(n859) );
  XNOR2_X1 U960 ( .A(KEYINPUT113), .B(n859), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U962 ( .A(KEYINPUT114), .B(n862), .Z(n928) );
  XNOR2_X1 U963 ( .A(n928), .B(n863), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(n921), .ZN(n868) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n866) );
  XNOR2_X1 U966 ( .A(G162), .B(KEYINPUT115), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n868), .B(n867), .Z(n871) );
  XOR2_X1 U969 ( .A(G164), .B(n869), .Z(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(n887) );
  NAND2_X1 U971 ( .A1(G118), .A2(n872), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G130), .A2(n873), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n882) );
  NAND2_X1 U974 ( .A1(G142), .A2(n876), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U977 ( .A(n880), .B(KEYINPUT45), .Z(n881) );
  NOR2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U980 ( .A(G160), .B(n885), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U982 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U983 ( .A(G301), .B(n889), .Z(n891) );
  XNOR2_X1 U984 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n892), .B(G286), .ZN(n893) );
  NOR2_X1 U986 ( .A1(G37), .A2(n893), .ZN(n894) );
  XNOR2_X1 U987 ( .A(KEYINPUT116), .B(n894), .ZN(G397) );
  XOR2_X1 U988 ( .A(G2438), .B(KEYINPUT108), .Z(n896) );
  XNOR2_X1 U989 ( .A(G1348), .B(G1341), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n906) );
  XOR2_X1 U991 ( .A(KEYINPUT110), .B(KEYINPUT107), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2446), .B(G2443), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U994 ( .A(G2430), .B(G2451), .Z(n900) );
  XNOR2_X1 U995 ( .A(G2454), .B(G2435), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U998 ( .A(KEYINPUT109), .B(G2427), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n907), .A2(G14), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(KEYINPUT117), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G96), .ZN(G221) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(n914), .ZN(G401) );
  INV_X1 U1013 ( .A(n915), .ZN(G223) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  INV_X1 U1015 ( .A(KEYINPUT55), .ZN(n941) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT51), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n938) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT118), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n936) );
  XOR2_X1 U1025 ( .A(G2072), .B(n928), .Z(n930) );
  XNOR2_X1 U1026 ( .A(G2078), .B(G164), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT50), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT119), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT52), .B(n939), .Z(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1036 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n955) );
  XOR2_X1 U1037 ( .A(G32), .B(G1996), .Z(n947) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(G27), .B(n943), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT120), .B(n950), .Z(n952) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n955), .B(n954), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G2084), .B(G34), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(KEYINPUT54), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(n961), .Z(n963) );
  INV_X1 U1055 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n964), .ZN(n1020) );
  INV_X1 U1058 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1059 ( .A(n1016), .B(KEYINPUT56), .Z(n990) );
  XOR2_X1 U1060 ( .A(n965), .B(G1341), .Z(n967) );
  XOR2_X1 U1061 ( .A(G301), .B(G1961), .Z(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n988) );
  XNOR2_X1 U1064 ( .A(G168), .B(G1966), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n972), .B(KEYINPUT122), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT57), .B(n973), .ZN(n983) );
  INV_X1 U1068 ( .A(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT123), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G1956), .B(G299), .Z(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n981) );
  XOR2_X1 U1073 ( .A(G1971), .B(G166), .Z(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1076 ( .A(G1348), .B(n984), .Z(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n1018) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1976), .B(G23), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n996), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT58), .ZN(n1010) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G21), .ZN(n1008) );
  XOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .Z(n998) );
  XNOR2_X1 U1090 ( .A(G4), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(G20), .B(G1956), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1006), .B(KEYINPUT124), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G5), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

