//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n439, new_n445, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  OR2_X1    g012(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(new_n439), .ZN(G220));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g016(.A(G69), .ZN(G235));
  INV_X1    g017(.A(G120), .ZN(G236));
  INV_X1    g018(.A(G57), .ZN(G237));
  XOR2_X1   g019(.A(KEYINPUT68), .B(G108), .Z(new_n445));
  INV_X1    g020(.A(new_n445), .ZN(G238));
  NAND4_X1  g021(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g029(.A1(G221), .A2(G218), .A3(G219), .ZN(new_n455));
  NAND3_X1  g030(.A1(new_n438), .A2(new_n455), .A3(new_n439), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  INV_X1    g038(.A(G567), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(new_n459), .ZN(new_n465));
  XOR2_X1   g040(.A(new_n465), .B(KEYINPUT70), .Z(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n474), .A2(new_n476), .A3(G137), .A4(new_n468), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n469), .A2(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n482), .A2(KEYINPUT71), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT71), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n474), .A2(new_n476), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n484), .A2(new_n485), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n474), .A2(new_n476), .A3(G126), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n474), .A2(new_n476), .A3(G138), .A4(new_n468), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n469), .A2(new_n501), .A3(G138), .A4(new_n468), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G651), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G543), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n506), .A2(new_n508), .B1(new_n505), .B2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G51), .A3(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(G89), .A3(new_n514), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n512), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n507), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n517), .A2(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT5), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n512), .A2(G43), .B1(G651), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n511), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n527), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT74), .B(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n544), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n517), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  NAND4_X1  g141(.A1(new_n509), .A2(G49), .A3(G543), .A4(new_n510), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n544), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n527), .A2(G48), .A3(G543), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n569), .ZN(G305));
  XOR2_X1   g155(.A(KEYINPUT76), .B(G47), .Z(new_n581));
  NAND2_X1  g156(.A1(new_n512), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n507), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n517), .A2(G85), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n569), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT77), .B(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n544), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G54), .B1(G651), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n587), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n587), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  XOR2_X1   g175(.A(G299), .B(KEYINPUT78), .Z(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  NAND2_X1  g178(.A1(new_n592), .A2(new_n596), .ZN(new_n604));
  INV_X1    g179(.A(G860), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(G559), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT79), .Z(G148));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n549), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n604), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n469), .A2(new_n478), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT13), .Z(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n487), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n486), .A2(G2105), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n468), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n617), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(G2100), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(G1341), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n634));
  INV_X1    g209(.A(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n633), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G14), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(KEYINPUT17), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n649), .ZN(new_n653));
  OAI21_X1  g228(.A(KEYINPUT18), .B1(new_n651), .B2(new_n648), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n648), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT83), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n671), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT21), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT22), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT84), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n676), .A2(new_n677), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n678), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n662), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n682), .B1(new_n679), .B2(new_n680), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n684), .A3(new_n678), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n661), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(G229));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G11), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT95), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(G28), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n694), .B2(G28), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n693), .B1(new_n695), .B2(new_n697), .C1(new_n622), .C2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n487), .A2(G129), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n478), .A2(G105), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT26), .ZN(new_n704));
  AOI211_X1 g279(.A(new_n702), .B(new_n704), .C1(G141), .C2(new_n618), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  OR2_X1    g283(.A1(G29), .A2(G32), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  AOI21_X1  g287(.A(new_n698), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  INV_X1    g289(.A(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G160), .B2(new_n696), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2084), .ZN(new_n719));
  INV_X1    g294(.A(new_n712), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n710), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n696), .A2(G27), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n500), .A2(new_n502), .ZN(new_n724));
  INV_X1    g299(.A(new_n498), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n723), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2078), .ZN(new_n728));
  NAND2_X1  g303(.A1(G168), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G21), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n713), .A2(new_n721), .A3(new_n728), .A4(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(G29), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n618), .A2(G139), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n478), .A2(G103), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n741), .A2(new_n742), .B1(new_n468), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n734), .B1(new_n744), .B2(new_n696), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2072), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n730), .A2(new_n731), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n597), .B2(new_n749), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT89), .B(G1348), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n733), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n550), .B2(new_n749), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1341), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n696), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n696), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n762), .A2(new_n763), .A3(G2090), .ZN(new_n764));
  OAI21_X1  g339(.A(G2090), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n696), .A2(G26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n618), .A2(G140), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n766), .B(new_n772), .S(KEYINPUT28), .Z(new_n773));
  XOR2_X1   g348(.A(KEYINPUT91), .B(G2067), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n749), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n749), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n764), .A2(new_n765), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n759), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT23), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n749), .A2(G20), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n782), .B(new_n783), .C1(G299), .C2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n782), .B2(new_n783), .ZN(new_n785));
  INV_X1    g360(.A(G1956), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n754), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n749), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n749), .ZN(new_n792));
  INV_X1    g367(.A(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G23), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT87), .Z(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n571), .B2(new_n749), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT33), .B(G1976), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n794), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n749), .A2(G24), .ZN(new_n806));
  INV_X1    g381(.A(G290), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n749), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT86), .B(G1986), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G25), .A2(G29), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n618), .A2(G131), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G119), .B2(new_n487), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n811), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT35), .B(G1991), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT85), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n808), .A2(new_n809), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n804), .A2(new_n805), .A3(new_n810), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT88), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n825), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n790), .B(KEYINPUT98), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n788), .B(KEYINPUT97), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n829), .B1(new_n826), .B2(new_n827), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(G311));
  OAI211_X1 g410(.A(new_n790), .B(KEYINPUT99), .C1(new_n828), .C2(new_n829), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(new_n597), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n544), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n512), .A2(G55), .B1(G651), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n517), .A2(G93), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n550), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n549), .A2(new_n847), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n851), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n605), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n771), .B(G164), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n706), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n744), .A2(KEYINPUT100), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n744), .A2(KEYINPUT100), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n816), .B(new_n614), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(G130), .A2(new_n487), .B1(new_n618), .B2(G142), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n468), .A2(KEYINPUT101), .A3(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n468), .B2(G118), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n622), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n491), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n865), .B2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g452(.A(G303), .B(G305), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n807), .A2(new_n571), .ZN(new_n880));
  INV_X1    g455(.A(new_n571), .ZN(new_n881));
  NAND2_X1  g456(.A1(G290), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(new_n882), .A3(new_n880), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n885), .A4(KEYINPUT42), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n849), .A2(new_n891), .A3(new_n850), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n849), .B2(new_n850), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n892), .A2(new_n893), .B1(G559), .B2(new_n604), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n851), .A2(KEYINPUT102), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n849), .A2(new_n891), .A3(new_n850), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n610), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n597), .A2(G299), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n604), .A2(new_n565), .A3(new_n561), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n894), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n894), .A2(new_n897), .A3(new_n904), .A4(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n894), .A2(new_n897), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n900), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n890), .A2(new_n907), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n905), .A2(new_n906), .B1(new_n909), .B2(new_n900), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  INV_X1    g489(.A(new_n890), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n890), .A4(new_n908), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(G868), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n848), .A2(new_n608), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(G295));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  AOI211_X1 g500(.A(KEYINPUT106), .B(new_n925), .C1(new_n919), .C2(G868), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(G331));
  NAND2_X1  g502(.A1(new_n884), .A2(new_n885), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G171), .A2(G286), .ZN(new_n930));
  NAND2_X1  g505(.A1(G168), .A2(G301), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n851), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n849), .A2(new_n850), .A3(new_n930), .A4(new_n931), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n902), .A2(new_n903), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n900), .A3(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n904), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n933), .A2(new_n900), .A3(new_n934), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n928), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n937), .A2(new_n941), .A3(new_n945), .A4(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(KEYINPUT107), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n949), .A3(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(KEYINPUT108), .A3(new_n946), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n943), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n948), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT109), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n953), .A2(new_n955), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n958), .B(new_n951), .C1(new_n959), .C2(new_n948), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(G397));
  INV_X1    g536(.A(KEYINPUT127), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n964));
  INV_X1    g539(.A(G125), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n471), .B1(new_n486), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G2105), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(G40), .A3(new_n479), .A4(new_n477), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n816), .B(new_n818), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n771), .B(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n707), .A2(G1996), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n706), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n974), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g554(.A(G290), .B(G1986), .Z(new_n980));
  AOI21_X1  g555(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT55), .ZN(new_n983));
  INV_X1    g558(.A(G40), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n472), .A2(new_n984), .A3(new_n480), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n964), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n726), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n793), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n726), .A2(new_n987), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n968), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n992));
  NOR3_X1   g567(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT112), .B(G2090), .Z(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n996), .A3(KEYINPUT116), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT116), .B1(new_n990), .B2(new_n996), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n983), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n990), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT111), .B(new_n793), .C1(new_n986), .C2(new_n989), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n996), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n983), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(G8), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G305), .A2(G1981), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n517), .A2(G86), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n578), .A4(new_n577), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n991), .A2(new_n968), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1007), .A2(new_n1010), .A3(KEYINPUT49), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n881), .A2(KEYINPUT113), .A3(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n724), .B2(new_n725), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n985), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n571), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1019), .A2(G8), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(G288), .A2(new_n1023), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1028), .A2(new_n1025), .A3(KEYINPUT52), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1000), .A2(new_n1006), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n968), .B1(new_n991), .B2(new_n963), .ZN(new_n1032));
  INV_X1    g607(.A(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n988), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n992), .A2(new_n994), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n778), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n988), .A2(KEYINPUT117), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1020), .A2(new_n1039), .A3(KEYINPUT45), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(new_n1038), .A3(new_n1033), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT125), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G301), .B(KEYINPUT54), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n1048));
  AND3_X1   g623(.A1(G286), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(G286), .B2(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n1051), .B2(KEYINPUT124), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n985), .B1(new_n1020), .B2(new_n1053), .ZN(new_n1054));
  OR3_X1    g629(.A1(new_n1054), .A2(G2084), .A3(new_n993), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1039), .B1(new_n1020), .B2(KEYINPUT45), .ZN(new_n1056));
  NOR4_X1   g631(.A1(G164), .A2(KEYINPUT117), .A3(new_n963), .A4(G1384), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n986), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1058), .B2(G1966), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1050), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G286), .A2(new_n1048), .A3(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1052), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1054), .A2(G2084), .A3(new_n993), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1032), .A2(new_n1040), .A3(new_n1038), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n731), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1051), .B1(new_n1066), .B2(new_n1015), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1051), .B(new_n1052), .C1(new_n1066), .C2(new_n1015), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1046), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1036), .A2(new_n778), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1033), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n468), .B1(new_n966), .B2(KEYINPUT126), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n480), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n964), .A3(new_n988), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1047), .A2(new_n1068), .A3(new_n1069), .A4(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n635), .B1(new_n1054), .B2(new_n993), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1014), .A2(new_n973), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n597), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1080), .A2(new_n1081), .A3(KEYINPUT60), .A4(new_n604), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1085), .B2(new_n597), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1084), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n786), .B1(new_n1054), .B2(new_n993), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(G2072), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n964), .A2(new_n988), .A3(new_n985), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n565), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G299), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n561), .B(new_n565), .C1(new_n1097), .C2(KEYINPUT57), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1102), .A2(new_n1104), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT121), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1103), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1106), .A2(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n964), .A2(new_n988), .A3(new_n976), .A4(new_n985), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(G1341), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1021), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n550), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT59), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1091), .A2(new_n1105), .A3(new_n1110), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1082), .A2(new_n597), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1108), .B1(new_n1119), .B2(new_n1102), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1079), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1062), .B1(new_n1059), .B2(G8), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1062), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1066), .B2(new_n1051), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT62), .B(new_n1069), .C1(new_n1123), .C2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1045), .A2(G171), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT62), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1031), .B1(new_n1122), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(G288), .B2(G1976), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(G288), .A2(new_n1135), .A3(G1976), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1010), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1016), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT114), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1142), .A2(new_n1019), .A3(new_n1024), .A4(new_n1016), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(new_n1026), .A4(new_n1018), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1146), .B2(new_n1006), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1004), .A2(G8), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1141), .B(new_n1145), .C1(new_n1148), .C2(new_n1005), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1066), .A2(new_n1015), .A3(G286), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1006), .A2(new_n1150), .A3(KEYINPUT63), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1000), .A2(new_n1006), .A3(new_n1030), .A4(new_n1150), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1147), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n981), .B1(new_n1133), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n969), .A2(new_n1159), .A3(KEYINPUT48), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT48), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1159), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n970), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1160), .B(new_n1163), .C1(new_n979), .C2(new_n970), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT46), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n970), .B2(G1996), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n969), .A2(KEYINPUT46), .A3(new_n976), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n707), .A2(new_n974), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1166), .B(new_n1167), .C1(new_n1168), .C2(new_n970), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT47), .ZN(new_n1170));
  INV_X1    g745(.A(new_n818), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n816), .A2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n978), .A2(new_n1172), .B1(G2067), .B2(new_n771), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n969), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1164), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n962), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1175), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1147), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(new_n1152), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1110), .A2(new_n1117), .A3(new_n1105), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1120), .B1(new_n1181), .B2(new_n1091), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n1182), .A2(new_n1079), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1180), .B1(new_n1183), .B2(new_n1031), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n1177), .C1(new_n1184), .C2(new_n981), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1176), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g761(.A(new_n466), .B(G227), .C1(new_n641), .C2(new_n643), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n687), .A2(new_n690), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n874), .B2(new_n875), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n1190), .A2(new_n950), .A3(new_n947), .ZN(G225));
  INV_X1    g765(.A(G225), .ZN(G308));
endmodule


