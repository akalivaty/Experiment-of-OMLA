//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n206), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT1), .B2(new_n203), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(KEYINPUT23), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n224));
  OR2_X1    g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(G176gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n216), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n235));
  OR2_X1    g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n233), .A2(new_n235), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n239), .B2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n237), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(new_n234), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n216), .A2(G176gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n226), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n241), .A2(new_n242), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT27), .B(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT28), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT28), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n220), .A2(KEYINPUT26), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n220), .A2(KEYINPUT26), .ZN(new_n257));
  INV_X1    g056(.A(new_n221), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n256), .B(new_n230), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n254), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n214), .B1(new_n249), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G227gat), .ZN(new_n262));
  INV_X1    g061(.A(G233gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n226), .B1(new_n228), .B2(new_n216), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n243), .A2(new_n232), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n266), .A2(KEYINPUT66), .B1(new_n267), .B2(new_n235), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT25), .B1(new_n268), .B2(new_n229), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n247), .B1(new_n269), .B2(KEYINPUT67), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n213), .B(new_n265), .C1(new_n270), .C2(new_n241), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n261), .A2(new_n264), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G15gat), .B(G43gat), .Z(new_n276));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n271), .ZN(new_n280));
  INV_X1    g079(.A(new_n264), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT34), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n264), .B1(new_n261), .B2(new_n271), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n278), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n272), .B(KEYINPUT32), .C1(new_n274), .C2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n279), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n279), .B2(new_n290), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT36), .ZN(new_n293));
  NOR3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n290), .ZN(new_n295));
  INV_X1    g094(.A(new_n288), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n288), .A3(new_n290), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT36), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(KEYINPUT2), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G141gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT72), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n307), .A2(KEYINPUT72), .A3(G141gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n300), .ZN(new_n312));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G141gat), .B(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT73), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT3), .A4(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n311), .A2(new_n320), .A3(new_n316), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n311), .B2(new_n316), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n311), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT74), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n322), .B(new_n213), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n210), .A2(new_n311), .A3(new_n316), .A4(new_n212), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n321), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n335), .B2(new_n214), .ZN(new_n336));
  INV_X1    g135(.A(new_n330), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n329), .A2(new_n334), .A3(new_n330), .A4(new_n332), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(KEYINPUT75), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n342), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT0), .ZN(new_n346));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n348), .A3(new_n343), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n352), .A2(new_n351), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n239), .A2(new_n240), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n248), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n260), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n365));
  XNOR2_X1  g164(.A(G197gat), .B(G204gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n265), .B1(new_n270), .B2(new_n241), .ZN(new_n374));
  INV_X1    g173(.A(new_n359), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n365), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n365), .B2(new_n376), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n358), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n359), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n373), .A3(new_n376), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n357), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n388), .A3(new_n357), .A4(new_n385), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n353), .A2(new_n354), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT31), .B(G50gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT3), .B1(new_n373), .B2(new_n381), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(new_n327), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n327), .B2(new_n325), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n373), .ZN(new_n398));
  INV_X1    g197(.A(G228gat), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n396), .A2(new_n398), .B1(new_n399), .B2(new_n263), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n263), .ZN(new_n401));
  OAI221_X1 g200(.A(new_n401), .B1(new_n397), .B2(new_n373), .C1(new_n335), .C2(new_n395), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT76), .B(G22gat), .Z(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n402), .ZN(new_n407));
  INV_X1    g206(.A(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n405), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n394), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n394), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(G22gat), .B2(new_n407), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI22_X1  g214(.A1(new_n294), .A2(new_n299), .B1(new_n390), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n353), .A2(new_n354), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n387), .A2(new_n389), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n415), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n293), .B1(new_n291), .B2(new_n292), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n297), .A2(KEYINPUT36), .A3(new_n298), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n426), .A3(KEYINPUT78), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n387), .A2(new_n389), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT79), .B(KEYINPUT39), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI211_X1 g231(.A(new_n330), .B(new_n432), .C1(new_n329), .C2(new_n332), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n433), .B2(new_n348), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n329), .A2(new_n332), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n337), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT80), .A3(new_n349), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n337), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n336), .A2(new_n337), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(KEYINPUT39), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n434), .A2(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n429), .B1(new_n441), .B2(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n438), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n433), .A2(new_n430), .A3(new_n348), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT80), .B1(new_n436), .B2(new_n349), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT40), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT81), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n341), .A2(KEYINPUT82), .A3(new_n343), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT82), .B1(new_n341), .B2(new_n343), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n348), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n441), .A2(KEYINPUT40), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n428), .A2(new_n449), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT37), .B1(new_n377), .B2(new_n378), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n384), .A2(new_n456), .A3(new_n385), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n358), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(new_n344), .B2(new_n349), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n455), .A2(new_n358), .A3(new_n457), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT38), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n463), .A2(new_n465), .A3(new_n354), .A4(new_n386), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n454), .B(new_n415), .C1(new_n461), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n418), .A2(new_n427), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n463), .A2(new_n354), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n412), .B2(new_n414), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n389), .B2(new_n387), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n297), .A2(KEYINPUT84), .A3(new_n298), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n291), .B2(new_n292), .ZN(new_n475));
  AND4_X1   g274(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n415), .A2(new_n297), .A3(new_n298), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT35), .B1(new_n421), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(KEYINPUT35), .C1(new_n421), .C2(new_n477), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n202), .B1(new_n468), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n481), .ZN(new_n484));
  INV_X1    g283(.A(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n418), .A2(new_n467), .A3(new_n427), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT86), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT88), .B(G29gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(G29gat), .A2(G36gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n491), .A2(new_n498), .A3(new_n496), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n493), .B(KEYINPUT89), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT17), .ZN(new_n502));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT7), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n505));
  XNOR2_X1  g304(.A(G99gat), .B(G106gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507));
  INV_X1    g306(.A(G85gat), .ZN(new_n508));
  INV_X1    g307(.A(G92gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(KEYINPUT8), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n510), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT96), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n502), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n511), .ZN(new_n516));
  AND2_X1   g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n516), .A2(new_n501), .B1(KEYINPUT41), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT97), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n517), .A2(KEYINPUT41), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT95), .ZN(new_n524));
  XOR2_X1   g323(.A(G134gat), .B(G162gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n519), .B(new_n520), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT93), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT16), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G1gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G1gat), .B2(new_n546), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G8gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n537), .B2(new_n536), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT94), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n529), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n536), .A2(new_n513), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n516), .B2(new_n536), .ZN(new_n561));
  INV_X1    g360(.A(G230gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n263), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n567));
  INV_X1    g366(.A(new_n536), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n514), .B2(new_n511), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(new_n560), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n516), .A2(KEYINPUT10), .A3(new_n568), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n566), .A2(new_n577), .A3(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n501), .A2(new_n550), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(new_n502), .B2(new_n551), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT90), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G113gat), .B(G141gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G197gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT11), .B(G169gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n501), .B(new_n550), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n588), .B(KEYINPUT13), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(KEYINPUT91), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n586), .A2(KEYINPUT18), .A3(new_n589), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n592), .A2(new_n598), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n590), .A2(new_n591), .B1(new_n604), .B2(new_n605), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(KEYINPUT92), .A3(new_n598), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(new_n598), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n583), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n489), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n419), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n428), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n624), .A2(G8gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G8gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT42), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(KEYINPUT42), .B2(new_n628), .ZN(G1325gat));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n426), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT100), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(G15gat), .B1(new_n619), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n475), .A2(new_n473), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n636), .A2(G15gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n619), .B2(new_n637), .ZN(G1326gat));
  NOR2_X1   g437(.A1(new_n619), .A2(new_n415), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT43), .B(G22gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1327gat));
  INV_X1    g440(.A(new_n492), .ZN(new_n642));
  INV_X1    g441(.A(new_n529), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n423), .A3(new_n467), .ZN(new_n644));
  AOI211_X1 g443(.A(KEYINPUT44), .B(new_n643), .C1(new_n486), .C2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n483), .A2(new_n488), .A3(new_n529), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(KEYINPUT44), .ZN(new_n647));
  INV_X1    g446(.A(new_n558), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(new_n617), .A3(new_n581), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n651), .B2(new_n621), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n489), .A2(new_n529), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n621), .A2(new_n642), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT45), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n653), .A2(KEYINPUT45), .A3(new_n654), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n655), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT101), .B1(new_n660), .B2(new_n652), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1328gat));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n650), .ZN(new_n663));
  INV_X1    g462(.A(G36gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n428), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT46), .Z(new_n666));
  NOR3_X1   g465(.A1(new_n647), .A2(new_n420), .A3(new_n650), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(G1329gat));
  INV_X1    g467(.A(new_n634), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n651), .A2(G43gat), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n636), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(G43gat), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g472(.A1(new_n651), .A2(new_n422), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G50gat), .ZN(new_n675));
  AOI211_X1 g474(.A(G50gat), .B(new_n415), .C1(new_n663), .C2(KEYINPUT102), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n663), .A2(KEYINPUT102), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(KEYINPUT103), .A2(KEYINPUT48), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT104), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(G1331gat));
  NAND2_X1  g485(.A1(new_n486), .A2(new_n644), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n617), .A2(new_n687), .A3(new_n559), .A4(new_n581), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n621), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g489(.A(new_n420), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n693), .B(new_n694), .Z(G1333gat));
  NAND2_X1  g494(.A1(new_n688), .A2(new_n669), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n636), .A2(G71gat), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n696), .A2(G71gat), .B1(new_n688), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g498(.A1(new_n688), .A2(new_n422), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT106), .B(G78gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1335gat));
  NAND2_X1  g501(.A1(new_n613), .A2(new_n616), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n648), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n581), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n706));
  INV_X1    g505(.A(new_n645), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n708), .B2(new_n621), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  NOR4_X1   g509(.A1(new_n647), .A2(new_n710), .A3(new_n419), .A4(new_n705), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n709), .A2(new_n711), .A3(new_n508), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n687), .A2(new_n529), .A3(new_n704), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n713), .A2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n714), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(KEYINPUT108), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n419), .A2(G85gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n717), .A2(new_n581), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT109), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n647), .A2(new_n419), .A3(new_n705), .ZN(new_n726));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726), .B2(KEYINPUT107), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n725), .B(new_n722), .C1(new_n727), .C2(new_n711), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1336gat));
  NAND4_X1  g528(.A1(new_n715), .A2(new_n509), .A3(new_n428), .A4(new_n581), .ZN(new_n730));
  INV_X1    g529(.A(new_n708), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n420), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(new_n509), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n730), .B2(KEYINPUT110), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI221_X1 g535(.A(new_n730), .B1(KEYINPUT110), .B2(new_n734), .C1(new_n732), .C2(new_n509), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1337gat));
  OAI21_X1  g537(.A(G99gat), .B1(new_n731), .B2(new_n634), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n717), .A2(new_n581), .A3(new_n720), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n636), .A2(G99gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(G1338gat));
  NAND2_X1  g541(.A1(new_n708), .A2(new_n422), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G106gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n582), .A2(G106gat), .A3(new_n415), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT53), .B1(new_n715), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n745), .B(KEYINPUT111), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n743), .A2(G106gat), .B1(new_n715), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(G1339gat));
  NOR2_X1   g550(.A1(new_n583), .A2(new_n703), .ZN(new_n752));
  INV_X1    g551(.A(new_n596), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n586), .A2(new_n589), .B1(new_n599), .B2(new_n601), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n610), .A2(new_n612), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n581), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n570), .A2(new_n563), .A3(new_n571), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n570), .A2(new_n759), .A3(new_n563), .A4(new_n571), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(new_n573), .A3(KEYINPUT54), .A4(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n577), .B1(new_n572), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n580), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n756), .B1(new_n769), .B2(new_n617), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n643), .ZN(new_n771));
  INV_X1    g570(.A(new_n769), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n529), .A3(new_n755), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n752), .B1(new_n774), .B2(new_n558), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n422), .ZN(new_n776));
  INV_X1    g575(.A(new_n636), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n428), .A2(new_n419), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G113gat), .B1(new_n779), .B2(new_n617), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n775), .A2(new_n419), .A3(new_n428), .A4(new_n477), .ZN(new_n781));
  INV_X1    g580(.A(G113gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n703), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT113), .ZN(G1340gat));
  NOR3_X1   g584(.A1(new_n779), .A2(new_n208), .A3(new_n582), .ZN(new_n786));
  AOI21_X1  g585(.A(G120gat), .B1(new_n781), .B2(new_n581), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(G1341gat));
  OAI21_X1  g587(.A(G127gat), .B1(new_n779), .B2(new_n558), .ZN(new_n789));
  INV_X1    g588(.A(G127gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n781), .A2(new_n790), .A3(new_n648), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1342gat));
  INV_X1    g591(.A(G134gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n781), .A2(new_n793), .A3(new_n529), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT114), .B(KEYINPUT56), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  OAI21_X1  g596(.A(G134gat), .B1(new_n779), .B2(new_n643), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(G1343gat));
  AOI21_X1  g598(.A(KEYINPUT55), .B1(new_n764), .B2(KEYINPUT115), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(KEYINPUT115), .B2(new_n764), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n703), .A3(new_n767), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n756), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n643), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n766), .B1(new_n616), .B2(new_n613), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n806), .A2(new_n801), .B1(new_n581), .B2(new_n755), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(KEYINPUT116), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n773), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n752), .B1(new_n809), .B2(new_n558), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n415), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n774), .A2(new_n558), .ZN(new_n815));
  INV_X1    g614(.A(new_n752), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT57), .B1(new_n817), .B2(new_n422), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n773), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n529), .B1(new_n807), .B2(KEYINPUT116), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n804), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n823), .B2(new_n648), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n812), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n814), .A2(new_n819), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n634), .A2(new_n778), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G141gat), .B1(new_n830), .B2(new_n617), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n669), .A2(new_n415), .ZN(new_n832));
  AND4_X1   g631(.A1(new_n621), .A2(new_n817), .A3(new_n420), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n305), .A3(new_n703), .ZN(new_n834));
  NAND2_X1  g633(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT119), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n836), .A3(new_n839), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1344gat));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n581), .A3(new_n829), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n307), .A2(KEYINPUT59), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n775), .A2(new_n813), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n824), .A2(new_n422), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n811), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n828), .A2(new_n582), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G148gat), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n845), .A2(new_n846), .B1(new_n852), .B2(KEYINPUT59), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n833), .A2(new_n307), .A3(new_n581), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n844), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n846), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n824), .A2(new_n812), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n818), .B1(KEYINPUT117), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n828), .B1(new_n859), .B2(new_n826), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n860), .B2(new_n581), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n811), .B1(new_n810), .B2(new_n415), .ZN(new_n863));
  INV_X1    g662(.A(new_n847), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n850), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n862), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n854), .C1(new_n861), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n856), .A2(new_n868), .ZN(G1345gat));
  OAI21_X1  g668(.A(G155gat), .B1(new_n830), .B2(new_n558), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n833), .A2(new_n301), .A3(new_n648), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1346gat));
  NAND3_X1  g671(.A1(new_n833), .A2(new_n302), .A3(new_n529), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n830), .A2(new_n643), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n875));
  OAI21_X1  g674(.A(G162gat), .B1(new_n874), .B2(KEYINPUT121), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n775), .A2(new_n621), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n477), .A2(new_n420), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(G169gat), .A3(new_n617), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n621), .A2(new_n420), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n777), .A2(KEYINPUT123), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885));
  INV_X1    g684(.A(new_n883), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n636), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n776), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n617), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT124), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n882), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1348gat));
  INV_X1    g693(.A(new_n880), .ZN(new_n895));
  AOI21_X1  g694(.A(G176gat), .B1(new_n895), .B2(new_n581), .ZN(new_n896));
  INV_X1    g695(.A(new_n888), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n581), .A2(new_n228), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1349gat));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n250), .A3(new_n648), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n888), .B2(new_n558), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n888), .B2(new_n643), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(KEYINPUT125), .B2(new_n904), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n880), .A2(G190gat), .A3(new_n643), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1351gat));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n669), .A2(new_n886), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n865), .A2(new_n703), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(KEYINPUT126), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(KEYINPUT126), .B2(new_n914), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n878), .A2(new_n428), .A3(new_n832), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n912), .A3(new_n703), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1352gat));
  INV_X1    g718(.A(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n920), .A3(new_n581), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT62), .Z(new_n922));
  NAND2_X1  g721(.A1(new_n865), .A2(new_n913), .ZN(new_n923));
  OAI21_X1  g722(.A(G204gat), .B1(new_n923), .B2(new_n582), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n368), .A3(new_n648), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n824), .B2(new_n422), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n648), .B(new_n913), .C1(new_n927), .C2(new_n847), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT127), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n923), .B2(new_n643), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n917), .A2(new_n369), .A3(new_n529), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


