//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n188), .A2(KEYINPUT68), .A3(new_n189), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n191), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n200), .A3(new_n202), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(G101), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G101), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n195), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  OR3_X1    g024(.A1(new_n210), .A2(KEYINPUT5), .A3(G119), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(KEYINPUT85), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(KEYINPUT85), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(G113), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT68), .B1(new_n188), .B2(new_n189), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n193), .A2(new_n187), .A3(new_n192), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n199), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n196), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(new_n203), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n203), .A2(new_n222), .A3(new_n219), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n215), .B(new_n218), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n209), .A2(new_n225), .A3(new_n227), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT65), .B(G143), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(G143), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT67), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT67), .A2(G128), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n238), .A2(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n235), .B2(G146), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n236), .A2(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G125), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT0), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n244), .A3(KEYINPUT64), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(KEYINPUT0), .B2(G128), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n251), .A2(new_n253), .B1(KEYINPUT0), .B2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n248), .B1(new_n256), .B2(new_n247), .ZN(new_n257));
  INV_X1    g071(.A(G224), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G953), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n257), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n226), .A2(new_n261), .A3(new_n228), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n231), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT7), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n248), .B(new_n265), .C1(new_n256), .C2(new_n247), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G143), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n270), .A3(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n237), .A3(new_n245), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n270), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n233), .B1(new_n273), .B2(new_n232), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n244), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT67), .A2(G128), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n276), .A2(new_n277), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n272), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G125), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n247), .B1(new_n249), .B2(new_n255), .ZN(new_n281));
  OAI22_X1  g095(.A1(new_n280), .A2(new_n281), .B1(new_n264), .B2(new_n259), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n230), .A2(new_n266), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n215), .A2(new_n218), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n203), .A2(new_n222), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n225), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n227), .B(KEYINPUT8), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n263), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G210), .B1(G237), .B2(G902), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n292), .B(KEYINPUT86), .Z(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G952), .ZN(new_n296));
  AOI211_X1 g110(.A(G953), .B(new_n296), .C1(G234), .C2(G237), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n298), .B(new_n299), .C1(G234), .C2(G237), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT21), .B(G898), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n263), .A2(new_n290), .A3(new_n293), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n295), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n307));
  INV_X1    g121(.A(G122), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n210), .A2(G122), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G107), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n309), .B(new_n310), .C1(KEYINPUT14), .C2(new_n199), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n268), .A2(new_n270), .A3(G128), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n276), .A2(G143), .A3(new_n277), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G134), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n315), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n240), .A2(new_n241), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n316), .A2(new_n323), .B1(new_n324), .B2(G143), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n235), .A2(KEYINPUT13), .A3(G128), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n309), .A2(new_n310), .A3(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n311), .A2(new_n199), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT92), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n316), .A2(new_n323), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n326), .A3(new_n317), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G134), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n328), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n322), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(G953), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n307), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n322), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n327), .A2(KEYINPUT92), .A3(new_n330), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n338), .B1(new_n334), .B2(new_n337), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n343), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n307), .A3(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n298), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT94), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT94), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n351), .A2(new_n355), .A3(new_n298), .A4(new_n352), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT15), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n354), .A2(new_n356), .B1(new_n357), .B2(G478), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT90), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n267), .A2(new_n361), .A3(new_n299), .A4(G214), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n235), .B2(KEYINPUT87), .ZN(new_n363));
  INV_X1    g177(.A(G214), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(G237), .A3(G953), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n235), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G131), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n363), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n365), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n273), .B2(KEYINPUT87), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n365), .B(new_n267), .C1(KEYINPUT65), .C2(new_n366), .ZN(new_n372));
  AOI21_X1  g186(.A(G131), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n360), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n247), .A2(G140), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT79), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n375), .A2(KEYINPUT79), .A3(G125), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT16), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n232), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G125), .B(G140), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n375), .A2(KEYINPUT79), .A3(G125), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n384), .B2(KEYINPUT79), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n389), .B2(new_n386), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n383), .B1(new_n232), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n368), .B1(new_n363), .B2(new_n367), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n371), .A2(G131), .A3(new_n372), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(KEYINPUT90), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n374), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n396), .B(new_n397), .C1(new_n363), .C2(new_n367), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n378), .A2(new_n379), .A3(G146), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(G146), .B2(new_n385), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n371), .A2(new_n372), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT18), .B(G131), .C1(new_n401), .C2(KEYINPUT88), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n403), .B(KEYINPUT89), .C1(new_n371), .C2(new_n372), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n398), .B(new_n400), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n196), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT91), .A4(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n380), .A2(new_n232), .A3(new_n382), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n383), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n392), .A2(new_n411), .A3(new_n393), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n408), .B(new_n405), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n359), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  AOI211_X1 g238(.A(KEYINPUT20), .B(new_n424), .C1(new_n410), .C2(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(G475), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n405), .B1(new_n416), .B2(new_n419), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n409), .ZN(new_n428));
  AOI21_X1  g242(.A(G902), .B1(new_n428), .B2(new_n420), .ZN(new_n429));
  OAI22_X1  g243(.A1(new_n423), .A2(new_n425), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n356), .A2(new_n357), .A3(G478), .ZN(new_n431));
  NOR4_X1   g245(.A1(new_n306), .A2(new_n358), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n204), .B(new_n207), .ZN(new_n434));
  INV_X1    g248(.A(new_n223), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n203), .A2(new_n222), .A3(new_n219), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT10), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n236), .A2(new_n242), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n272), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n434), .A2(new_n256), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT66), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n318), .A2(G137), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(KEYINPUT66), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT11), .A4(G134), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n318), .A2(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n446), .A2(new_n451), .A3(G131), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n448), .A2(G134), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n443), .B2(new_n444), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n447), .A2(KEYINPUT11), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n448), .A2(G134), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n368), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n271), .A2(new_n237), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n239), .B1(new_n273), .B2(new_n232), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n244), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n463), .A2(new_n464), .B1(new_n243), .B2(new_n245), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT80), .B(new_n461), .C1(new_n462), .C2(new_n244), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n285), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n441), .B(new_n460), .C1(new_n467), .C2(KEYINPUT10), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n299), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(KEYINPUT83), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n279), .A2(new_n224), .A3(new_n223), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n269), .A2(G143), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n232), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n244), .B1(new_n478), .B2(KEYINPUT1), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n464), .B1(new_n479), .B2(new_n243), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n272), .A3(new_n466), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n475), .B1(new_n481), .B2(new_n286), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n482), .B2(new_n460), .ZN(new_n483));
  INV_X1    g297(.A(new_n460), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT12), .B(new_n484), .C1(new_n467), .C2(new_n475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT83), .B1(new_n468), .B2(new_n472), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n433), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n472), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT84), .A3(new_n486), .A4(new_n473), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n441), .B1(new_n467), .B2(KEYINPUT10), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n468), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n471), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n298), .ZN(new_n500));
  NAND2_X1  g314(.A1(G469), .A2(G902), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n486), .A2(new_n502), .A3(new_n468), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n486), .B2(new_n468), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n471), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n490), .B1(new_n484), .B2(new_n494), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(G469), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n501), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G221), .ZN(new_n511));
  INV_X1    g325(.A(new_n341), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n298), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n432), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n342), .B1(G234), .B2(new_n298), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n383), .B1(new_n232), .B2(new_n384), .ZN(new_n517));
  INV_X1    g331(.A(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G128), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(G128), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n324), .A2(G119), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT23), .ZN(new_n523));
  OAI221_X1 g337(.A(new_n519), .B1(new_n520), .B2(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G110), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT24), .B(G110), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT77), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(KEYINPUT76), .A3(G128), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n522), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n324), .A2(KEYINPUT75), .A3(G119), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n524), .A2(G110), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n527), .A3(new_n533), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n413), .C2(new_n383), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT22), .B(G137), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n540), .B(new_n541), .Z(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n535), .B2(new_n538), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT25), .B1(new_n546), .B2(new_n298), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NOR4_X1   g362(.A1(new_n544), .A2(new_n545), .A3(new_n548), .A4(G902), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n516), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n516), .A2(G902), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n195), .A2(KEYINPUT70), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n249), .B(new_n255), .C1(new_n452), .C2(new_n459), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n454), .A2(new_n368), .A3(new_n458), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n444), .B2(new_n453), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n279), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n218), .A2(new_n559), .A3(new_n190), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n554), .A2(new_n555), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n558), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n561), .A2(new_n562), .B1(new_n195), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n279), .A2(KEYINPUT69), .A3(new_n556), .A4(new_n557), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n555), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n556), .A2(new_n557), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT69), .B1(new_n567), .B2(new_n279), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n554), .A2(new_n560), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n564), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n361), .A2(new_n299), .A3(G210), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT27), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n195), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT30), .B1(new_n566), .B2(new_n568), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT30), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n555), .A2(new_n558), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n580), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n556), .A2(new_n557), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n246), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n565), .A3(new_n555), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n570), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n584), .A2(new_n589), .A3(new_n578), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n579), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n581), .A2(new_n583), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n593), .B2(new_n195), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n591), .A4(new_n577), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n555), .A2(new_n558), .A3(new_n582), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(KEYINPUT30), .B2(new_n588), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n572), .B(new_n577), .C1(new_n598), .C2(new_n580), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT71), .B1(new_n599), .B2(KEYINPUT31), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n592), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(G472), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT32), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n600), .A2(new_n596), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n599), .A2(KEYINPUT31), .B1(new_n573), .B2(new_n578), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT32), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n588), .A2(new_n570), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n572), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT28), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n561), .A2(KEYINPUT73), .A3(new_n562), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT73), .B1(new_n561), .B2(new_n562), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT29), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n578), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n619), .B2(KEYINPUT74), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n578), .B1(new_n584), .B2(new_n589), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n564), .B(new_n577), .C1(new_n572), .C2(new_n562), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT72), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT74), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n613), .A2(new_n625), .A3(new_n616), .A4(new_n618), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT72), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n621), .A2(new_n627), .A3(new_n622), .A4(new_n617), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n620), .A2(new_n624), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n553), .B1(new_n610), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n515), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NAND2_X1  g447(.A1(new_n510), .A2(new_n514), .ZN(new_n634));
  INV_X1    g448(.A(new_n607), .ZN(new_n635));
  INV_X1    g449(.A(new_n553), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n605), .B2(new_n606), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT95), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(G128), .B1(new_n237), .B2(new_n271), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n272), .B1(new_n642), .B2(KEYINPUT80), .ZN(new_n643));
  INV_X1    g457(.A(new_n466), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n286), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n475), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT12), .B1(new_n647), .B2(new_n484), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n482), .A2(new_n474), .A3(new_n460), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n468), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT82), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n503), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n507), .B1(new_n652), .B2(new_n471), .ZN(new_n653));
  OAI21_X1  g467(.A(G469), .B1(new_n653), .B2(G902), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n513), .B1(new_n654), .B2(new_n500), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n605), .A2(new_n606), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n637), .B1(new_n656), .B2(new_n298), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n607), .A3(new_n553), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n351), .A2(new_n662), .A3(new_n352), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n345), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n340), .A2(KEYINPUT97), .A3(new_n343), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT96), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n348), .B2(new_n349), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n340), .A2(KEYINPUT96), .A3(new_n343), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n666), .B(new_n667), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(G478), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n663), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n353), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n430), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n306), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n661), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT34), .B(G104), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  INV_X1    g495(.A(new_n430), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n358), .B2(new_n431), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n306), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n661), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT35), .B(G107), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  NOR2_X1   g501(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n539), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n551), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n550), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n657), .A2(new_n692), .A3(new_n607), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n515), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT37), .B(G110), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G12));
  AOI21_X1  g511(.A(new_n608), .B1(new_n656), .B2(new_n602), .ZN(new_n698));
  AOI211_X1 g512(.A(KEYINPUT32), .B(new_n603), .C1(new_n605), .C2(new_n606), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n630), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n297), .B1(new_n300), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n682), .B(new_n703), .C1(new_n358), .C2(new_n431), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n295), .A2(new_n305), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n691), .A2(new_n706), .A3(new_n304), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n655), .A2(new_n700), .A3(new_n705), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XOR2_X1   g524(.A(new_n702), .B(KEYINPUT39), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n655), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n612), .A2(new_n578), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n599), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n717));
  AOI21_X1  g531(.A(G902), .B1(new_n716), .B2(KEYINPUT99), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI22_X1  g533(.A1(new_n698), .A2(new_n699), .B1(new_n637), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n706), .B(KEYINPUT38), .Z(new_n721));
  INV_X1    g535(.A(new_n304), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n430), .B1(new_n358), .B2(new_n431), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n691), .A4(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n713), .A2(new_n714), .A3(new_n720), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n273), .ZN(G45));
  INV_X1    g540(.A(KEYINPUT100), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n408), .B1(new_n395), .B2(new_n405), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n398), .A2(new_n400), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n363), .A2(new_n367), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n397), .B1(new_n730), .B2(new_n403), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n401), .A2(KEYINPUT88), .A3(new_n396), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n417), .A2(new_n418), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n728), .B1(new_n736), .B2(new_n408), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT20), .B1(new_n737), .B2(new_n424), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n421), .A2(new_n359), .A3(new_n422), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n428), .A2(new_n420), .ZN(new_n741));
  OAI21_X1  g555(.A(G475), .B1(new_n741), .B2(G902), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n740), .A2(new_n742), .B1(new_n674), .B2(new_n675), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n727), .B1(new_n743), .B2(new_n703), .ZN(new_n744));
  AND4_X1   g558(.A1(new_n727), .A2(new_n676), .A3(new_n430), .A4(new_n703), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n655), .A2(new_n746), .A3(new_n700), .A4(new_n708), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  NAND2_X1  g562(.A1(KEYINPUT101), .A2(G469), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n498), .A2(new_n298), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n749), .B1(new_n498), .B2(new_n298), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n751), .A3(new_n513), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n700), .A3(new_n636), .A4(new_n678), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n700), .A3(new_n684), .A4(new_n636), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  OR2_X1    g571(.A1(new_n358), .A2(new_n431), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n302), .A3(new_n430), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n759), .A3(new_n700), .A4(new_n708), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G119), .ZN(G21));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n602), .B(KEYINPUT102), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n613), .A2(new_n616), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n765), .A2(new_n578), .B1(KEYINPUT31), .B2(new_n599), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n766), .B2(new_n605), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n656), .A2(new_n298), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(G472), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT103), .B1(new_n769), .B2(new_n636), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n657), .A2(new_n767), .A3(new_n771), .A4(new_n553), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n723), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT104), .B(new_n430), .C1(new_n358), .C2(new_n431), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n302), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n706), .A2(new_n304), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(new_n752), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n762), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n767), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n771), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n769), .A2(KEYINPUT103), .A3(new_n636), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n752), .A2(new_n779), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n777), .A4(KEYINPUT105), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  NOR3_X1   g604(.A1(new_n657), .A2(new_n692), .A3(new_n767), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n752), .A2(new_n746), .A3(new_n791), .A4(new_n779), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G125), .ZN(G27));
  NOR2_X1   g607(.A1(new_n706), .A2(new_n722), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n700), .A2(new_n636), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT42), .A3(new_n655), .A4(new_n746), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT42), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n655), .A2(new_n700), .A3(new_n636), .A4(new_n794), .ZN(new_n798));
  INV_X1    g612(.A(new_n746), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  INV_X1    g616(.A(new_n798), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n704), .B(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  OR2_X1    g620(.A1(new_n653), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n653), .A2(KEYINPUT45), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(G469), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT46), .B1(new_n809), .B2(new_n501), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT107), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(KEYINPUT46), .A3(new_n501), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n500), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n514), .ZN(new_n816));
  INV_X1    g630(.A(new_n711), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n816), .A2(KEYINPUT108), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT108), .B1(new_n816), .B2(new_n817), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n430), .B1(new_n675), .B2(new_n674), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT43), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n430), .B2(KEYINPUT109), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n820), .B(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n823), .B(new_n691), .C1(new_n607), .C2(new_n657), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT44), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n794), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(new_n819), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G137), .ZN(G39));
  INV_X1    g644(.A(KEYINPUT47), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n816), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n514), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n794), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n799), .A2(new_n700), .A3(new_n636), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n752), .A2(new_n794), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT115), .ZN(new_n841));
  INV_X1    g655(.A(new_n297), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n840), .B2(KEYINPUT115), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n791), .A3(new_n823), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n786), .A2(new_n297), .A3(new_n823), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n722), .A3(new_n721), .A4(new_n752), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n845), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n720), .A2(new_n553), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n676), .A2(new_n430), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n841), .A2(new_n843), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT116), .Z(new_n858));
  OAI21_X1  g672(.A(new_n839), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n853), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n851), .ZN(new_n861));
  INV_X1    g675(.A(new_n858), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n862), .A4(new_n845), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  OR3_X1    g678(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT113), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT113), .B1(new_n750), .B2(new_n751), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n513), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n832), .A2(new_n833), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n847), .A2(new_n794), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n859), .A2(new_n863), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n844), .A2(new_n631), .A3(new_n823), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n876), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n844), .A2(new_n743), .A3(new_n855), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n296), .B(G953), .C1(new_n847), .C2(new_n787), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n868), .A2(new_n870), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n862), .A3(new_n861), .A4(new_n845), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n883), .B2(new_n864), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n778), .B1(new_n775), .B2(new_n776), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n691), .A2(new_n702), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n655), .A3(new_n720), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n792), .A3(new_n747), .A4(new_n709), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n758), .A2(new_n430), .A3(new_n702), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n700), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n746), .A2(new_n769), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n634), .A2(new_n692), .A3(new_n835), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n803), .A2(new_n804), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n890), .A2(new_n801), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT111), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n678), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n677), .A2(new_n306), .A3(KEYINPUT111), .ZN(new_n900));
  OAI22_X1  g714(.A1(new_n899), .A2(new_n900), .B1(new_n306), .B2(new_n683), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n640), .A2(new_n660), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n631), .B(new_n752), .C1(new_n678), .C2(new_n684), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n515), .B1(new_n631), .B2(new_n693), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n760), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n781), .B2(new_n788), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n707), .B1(new_n610), .B2(new_n630), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(new_n655), .C1(new_n705), .C2(new_n746), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n792), .A4(new_n888), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n897), .A2(new_n906), .A3(KEYINPUT53), .A4(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n890), .A2(new_n801), .A3(new_n896), .A4(new_n910), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n760), .A2(new_n753), .A3(new_n756), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n655), .A2(new_n432), .ZN(new_n915));
  INV_X1    g729(.A(new_n693), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n700), .A2(new_n636), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n789), .A2(new_n919), .A3(new_n902), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n912), .B1(new_n913), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n911), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n923), .B(new_n925), .C1(new_n872), .C2(KEYINPUT118), .ZN(new_n926));
  OAI22_X1  g740(.A1(new_n885), .A2(new_n926), .B1(G952), .B2(G953), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n750), .A2(new_n751), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT49), .Z(new_n929));
  NAND4_X1  g743(.A1(new_n636), .A2(new_n820), .A3(new_n514), .A4(new_n304), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT110), .Z(new_n931));
  INV_X1    g745(.A(new_n721), .ZN(new_n932));
  OR4_X1    g746(.A1(new_n720), .A2(new_n929), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n933), .ZN(G75));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n922), .A2(G902), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n294), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n231), .A2(new_n262), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n260), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT55), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n937), .A2(new_n940), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n299), .A2(G952), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G51));
  INV_X1    g758(.A(new_n924), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n922), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n501), .B(KEYINPUT57), .Z(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n498), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n936), .A2(new_n809), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(G54));
  NAND4_X1  g768(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n737), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n737), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n943), .ZN(G60));
  AND2_X1   g772(.A1(new_n663), .A2(new_n671), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n947), .A2(new_n949), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n943), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n923), .B2(new_n925), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n959), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT121), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n967), .A2(new_n959), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT121), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(new_n971), .A3(new_n966), .A4(new_n964), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n911), .B2(new_n921), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n689), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT61), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n966), .B1(new_n978), .B2(new_n546), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n981), .A2(KEYINPUT123), .B1(new_n689), .B2(new_n978), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n985), .B(new_n966), .C1(new_n978), .C2(new_n546), .ZN(new_n986));
  AOI211_X1 g800(.A(new_n983), .B(KEYINPUT61), .C1(new_n984), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n981), .A2(KEYINPUT123), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n986), .A3(new_n979), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT124), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n982), .B1(new_n987), .B2(new_n991), .ZN(G66));
  OAI21_X1  g806(.A(G953), .B1(new_n301), .B2(new_n258), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT125), .Z(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n920), .B2(new_n299), .ZN(new_n995));
  INV_X1    g809(.A(G898), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n938), .B1(new_n996), .B2(G953), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G69));
  AND2_X1   g812(.A1(new_n908), .A2(new_n792), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n725), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT62), .Z(new_n1001));
  AOI21_X1  g815(.A(new_n743), .B1(new_n758), .B2(new_n682), .ZN(new_n1002));
  OR4_X1    g816(.A1(new_n917), .A2(new_n712), .A3(new_n835), .A4(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n829), .A2(new_n837), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n299), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n598), .B(new_n390), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(G900), .B2(G953), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n999), .A2(new_n801), .A3(new_n805), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n818), .A2(new_n819), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n828), .B1(new_n631), .B2(new_n886), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n837), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1008), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n299), .B1(G227), .B2(G900), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1015), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1007), .A2(new_n1017), .A3(new_n1013), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(new_n594), .A2(new_n578), .ZN(new_n1020));
  XNOR2_X1  g834(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n637), .A2(new_n298), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1012), .B2(new_n920), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g841(.A(KEYINPUT127), .B(new_n1024), .C1(new_n1012), .C2(new_n920), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1024), .B1(new_n1004), .B2(new_n920), .ZN(new_n1030));
  INV_X1    g844(.A(new_n594), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1030), .A2(new_n1031), .A3(new_n577), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1023), .B1(new_n621), .B2(new_n599), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n943), .B1(new_n922), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1029), .A2(new_n1035), .ZN(G57));
endmodule


