

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  INV_X1 U328 ( .A(G204GAT), .ZN(n362) );
  XNOR2_X1 U329 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U330 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U331 ( .A(n369), .B(KEYINPUT26), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n371), .B(n370), .ZN(n572) );
  NOR2_X1 U333 ( .A1(n501), .A2(n470), .ZN(n463) );
  XNOR2_X1 U334 ( .A(KEYINPUT108), .B(G36GAT), .ZN(n464) );
  XNOR2_X1 U335 ( .A(n465), .B(n464), .ZN(G1329GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n297) );
  XNOR2_X1 U337 ( .A(KEYINPUT18), .B(G169GAT), .ZN(n296) );
  XNOR2_X1 U338 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U339 ( .A(KEYINPUT17), .B(n298), .Z(n324) );
  XOR2_X1 U340 ( .A(KEYINPUT21), .B(G197GAT), .Z(n354) );
  XOR2_X1 U341 ( .A(KEYINPUT94), .B(n354), .Z(n300) );
  NAND2_X1 U342 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U344 ( .A(KEYINPUT74), .B(G204GAT), .Z(n302) );
  XNOR2_X1 U345 ( .A(G92GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U347 ( .A(G64GAT), .B(n303), .Z(n438) );
  XOR2_X1 U348 ( .A(n304), .B(n438), .Z(n308) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(G36GAT), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n305), .B(G190GAT), .ZN(n414) );
  XNOR2_X1 U351 ( .A(G183GAT), .B(G211GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n306), .B(G8GAT), .ZN(n391) );
  XNOR2_X1 U353 ( .A(n414), .B(n391), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n324), .B(n309), .ZN(n548) );
  XOR2_X1 U356 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n311) );
  XNOR2_X1 U357 ( .A(G190GAT), .B(G71GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(G127GAT), .B(G15GAT), .Z(n390) );
  XOR2_X1 U360 ( .A(n312), .B(n390), .Z(n314) );
  XNOR2_X1 U361 ( .A(G43GAT), .B(G99GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U363 ( .A(G113GAT), .B(G120GAT), .Z(n316) );
  XNOR2_X1 U364 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n336) );
  XOR2_X1 U366 ( .A(n336), .B(G176GAT), .Z(n318) );
  NAND2_X1 U367 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(n320), .B(n319), .Z(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n322) );
  XNOR2_X1 U371 ( .A(G183GAT), .B(KEYINPUT64), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n557) );
  XOR2_X1 U375 ( .A(G1GAT), .B(KEYINPUT5), .Z(n328) );
  XNOR2_X1 U376 ( .A(G155GAT), .B(G148GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U378 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n330) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n343) );
  XNOR2_X1 U382 ( .A(G127GAT), .B(G29GAT), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n333), .B(G162GAT), .ZN(n335) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n334), .B(KEYINPUT2), .ZN(n361) );
  XOR2_X1 U386 ( .A(n335), .B(n361), .Z(n341) );
  XOR2_X1 U387 ( .A(n336), .B(KEYINPUT1), .Z(n338) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n339), .B(G85GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n554) );
  XNOR2_X1 U393 ( .A(KEYINPUT27), .B(n548), .ZN(n372) );
  NAND2_X1 U394 ( .A1(n554), .A2(n372), .ZN(n344) );
  XNOR2_X1 U395 ( .A(KEYINPUT95), .B(n344), .ZN(n533) );
  XOR2_X1 U396 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n346) );
  XNOR2_X1 U397 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n367) );
  XNOR2_X1 U399 ( .A(G148GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n347), .B(KEYINPUT73), .ZN(n434) );
  INV_X1 U401 ( .A(n434), .ZN(n348) );
  XOR2_X1 U402 ( .A(G162GAT), .B(G50GAT), .Z(n410) );
  NAND2_X1 U403 ( .A1(n348), .A2(n410), .ZN(n351) );
  INV_X1 U404 ( .A(n410), .ZN(n349) );
  NAND2_X1 U405 ( .A1(n434), .A2(n349), .ZN(n350) );
  NAND2_X1 U406 ( .A1(n351), .A2(n350), .ZN(n353) );
  NAND2_X1 U407 ( .A1(G228GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n356) );
  XOR2_X1 U410 ( .A(G155GAT), .B(G22GAT), .Z(n394) );
  XNOR2_X1 U411 ( .A(n394), .B(n354), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U414 ( .A(G218GAT), .B(G211GAT), .Z(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n361), .B(G78GAT), .ZN(n363) );
  XOR2_X1 U417 ( .A(n367), .B(n366), .Z(n555) );
  XNOR2_X1 U418 ( .A(n555), .B(KEYINPUT28), .ZN(n476) );
  NAND2_X1 U419 ( .A1(n533), .A2(n476), .ZN(n523) );
  NOR2_X1 U420 ( .A1(n557), .A2(n523), .ZN(n368) );
  XOR2_X1 U421 ( .A(KEYINPUT96), .B(n368), .Z(n383) );
  NOR2_X1 U422 ( .A1(n557), .A2(n555), .ZN(n371) );
  INV_X1 U423 ( .A(KEYINPUT97), .ZN(n369) );
  INV_X1 U424 ( .A(n554), .ZN(n378) );
  AND2_X1 U425 ( .A1(n372), .A2(n378), .ZN(n373) );
  NAND2_X1 U426 ( .A1(n572), .A2(n373), .ZN(n380) );
  NAND2_X1 U427 ( .A1(n548), .A2(n557), .ZN(n374) );
  NAND2_X1 U428 ( .A1(n374), .A2(n555), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n375), .B(KEYINPUT98), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n376), .B(KEYINPUT25), .ZN(n377) );
  NAND2_X1 U431 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U432 ( .A1(n380), .A2(n379), .ZN(n381) );
  XNOR2_X1 U433 ( .A(n381), .B(KEYINPUT99), .ZN(n382) );
  NAND2_X1 U434 ( .A1(n383), .A2(n382), .ZN(n384) );
  XNOR2_X1 U435 ( .A(KEYINPUT100), .B(n384), .ZN(n467) );
  XOR2_X1 U436 ( .A(KEYINPUT12), .B(KEYINPUT85), .Z(n386) );
  XNOR2_X1 U437 ( .A(KEYINPUT84), .B(KEYINPUT82), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n399) );
  XOR2_X1 U439 ( .A(KEYINPUT83), .B(KEYINPUT14), .Z(n388) );
  XNOR2_X1 U440 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U442 ( .A(G1GAT), .B(KEYINPUT69), .Z(n454) );
  XOR2_X1 U443 ( .A(n389), .B(n454), .Z(n397) );
  XOR2_X1 U444 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U445 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U449 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U450 ( .A(G78GAT), .B(G71GAT), .Z(n401) );
  XNOR2_X1 U451 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U453 ( .A(G57GAT), .B(n402), .ZN(n441) );
  XOR2_X1 U454 ( .A(n403), .B(n441), .Z(n542) );
  INV_X1 U455 ( .A(n542), .ZN(n585) );
  NAND2_X1 U456 ( .A1(n467), .A2(n585), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n404), .B(KEYINPUT103), .ZN(n423) );
  XOR2_X1 U458 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n406) );
  XNOR2_X1 U459 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(n407), .ZN(n460) );
  XOR2_X1 U462 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT10), .B(KEYINPUT79), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n421) );
  XOR2_X1 U465 ( .A(G92GAT), .B(G106GAT), .Z(n412) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G99GAT), .Z(n433) );
  XNOR2_X1 U467 ( .A(n410), .B(n433), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(n413), .B(KEYINPUT80), .Z(n419) );
  XOR2_X1 U470 ( .A(n414), .B(KEYINPUT9), .Z(n416) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U473 ( .A(G134GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n460), .B(n422), .ZN(n568) );
  XOR2_X1 U477 ( .A(KEYINPUT36), .B(n568), .Z(n587) );
  NAND2_X1 U478 ( .A1(n423), .A2(n587), .ZN(n426) );
  XOR2_X1 U479 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT37), .B(n424), .ZN(n425) );
  XOR2_X1 U481 ( .A(n426), .B(n425), .Z(n501) );
  XOR2_X1 U482 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n428) );
  XNOR2_X1 U483 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U485 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n430) );
  XNOR2_X1 U486 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U488 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U489 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U490 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n578) );
  XOR2_X1 U495 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n444) );
  XNOR2_X1 U496 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n458) );
  XOR2_X1 U498 ( .A(G169GAT), .B(G15GAT), .Z(n446) );
  XNOR2_X1 U499 ( .A(G36GAT), .B(G50GAT), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U501 ( .A(G197GAT), .B(G22GAT), .Z(n448) );
  XNOR2_X1 U502 ( .A(G113GAT), .B(G141GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U504 ( .A(n450), .B(n449), .Z(n456) );
  XOR2_X1 U505 ( .A(KEYINPUT70), .B(KEYINPUT66), .Z(n452) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U510 ( .A(n458), .B(n457), .Z(n459) );
  XOR2_X1 U511 ( .A(n460), .B(n459), .Z(n535) );
  INV_X1 U512 ( .A(n535), .ZN(n574) );
  NOR2_X1 U513 ( .A1(n578), .A2(n574), .ZN(n461) );
  XOR2_X1 U514 ( .A(n461), .B(KEYINPUT78), .Z(n470) );
  XNOR2_X1 U515 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n462) );
  XNOR2_X2 U516 ( .A(n463), .B(n462), .ZN(n486) );
  NAND2_X1 U517 ( .A1(n548), .A2(n486), .ZN(n465) );
  INV_X1 U518 ( .A(n568), .ZN(n544) );
  NOR2_X1 U519 ( .A1(n544), .A2(n585), .ZN(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT16), .B(n466), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U522 ( .A(n469), .B(KEYINPUT101), .Z(n488) );
  NOR2_X1 U523 ( .A1(n488), .A2(n470), .ZN(n477) );
  NAND2_X1 U524 ( .A1(n554), .A2(n477), .ZN(n471) );
  XNOR2_X1 U525 ( .A(KEYINPUT34), .B(n471), .ZN(n472) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(n472), .ZN(G1324GAT) );
  NAND2_X1 U527 ( .A1(n548), .A2(n477), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U529 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U530 ( .A1(n477), .A2(n557), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  INV_X1 U532 ( .A(n476), .ZN(n506) );
  NAND2_X1 U533 ( .A1(n477), .A2(n506), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(KEYINPUT107), .Z(n480) );
  XNOR2_X1 U536 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n486), .A2(n554), .ZN(n481) );
  XOR2_X1 U539 ( .A(n482), .B(n481), .Z(G1328GAT) );
  NAND2_X1 U540 ( .A1(n486), .A2(n557), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G43GAT), .B(n485), .ZN(G1330GAT) );
  NAND2_X1 U544 ( .A1(n486), .A2(n506), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U546 ( .A(n578), .B(KEYINPUT41), .ZN(n561) );
  INV_X1 U547 ( .A(n561), .ZN(n537) );
  NAND2_X1 U548 ( .A1(n574), .A2(n537), .ZN(n500) );
  NOR2_X1 U549 ( .A1(n500), .A2(n488), .ZN(n496) );
  NAND2_X1 U550 ( .A1(n496), .A2(n554), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT42), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1332GAT) );
  XOR2_X1 U554 ( .A(G64GAT), .B(KEYINPUT111), .Z(n493) );
  NAND2_X1 U555 ( .A1(n496), .A2(n548), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1333GAT) );
  NAND2_X1 U557 ( .A1(n496), .A2(n557), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT112), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G71GAT), .B(n495), .ZN(G1334GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n498) );
  NAND2_X1 U561 ( .A1(n496), .A2(n506), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U563 ( .A(G78GAT), .B(n499), .Z(G1335GAT) );
  NOR2_X1 U564 ( .A1(n501), .A2(n500), .ZN(n507) );
  NAND2_X1 U565 ( .A1(n507), .A2(n554), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U567 ( .A1(n548), .A2(n507), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n557), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT114), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G99GAT), .B(n505), .ZN(G1338GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n509) );
  NAND2_X1 U573 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G106GAT), .B(n510), .ZN(G1339GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT116), .B(n542), .Z(n565) );
  NAND2_X1 U577 ( .A1(n537), .A2(n535), .ZN(n511) );
  XOR2_X1 U578 ( .A(KEYINPUT46), .B(n511), .Z(n512) );
  NOR2_X1 U579 ( .A1(n544), .A2(n512), .ZN(n513) );
  NAND2_X1 U580 ( .A1(n565), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT47), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n587), .A2(n542), .ZN(n517) );
  XOR2_X1 U583 ( .A(KEYINPUT117), .B(KEYINPUT45), .Z(n515) );
  XNOR2_X1 U584 ( .A(KEYINPUT65), .B(n515), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U586 ( .A1(n518), .A2(n574), .ZN(n519) );
  NOR2_X1 U587 ( .A1(n519), .A2(n578), .ZN(n520) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT48), .B(n522), .ZN(n550) );
  NOR2_X1 U590 ( .A1(n523), .A2(n550), .ZN(n524) );
  NAND2_X1 U591 ( .A1(n557), .A2(n524), .ZN(n530) );
  NOR2_X1 U592 ( .A1(n574), .A2(n530), .ZN(n525) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n525), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n561), .A2(n530), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n565), .A2(n530), .ZN(n528) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(n528), .Z(n529) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  NOR2_X1 U600 ( .A1(n568), .A2(n530), .ZN(n532) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(G1343GAT) );
  NAND2_X1 U603 ( .A1(n533), .A2(n572), .ZN(n534) );
  NOR2_X1 U604 ( .A1(n550), .A2(n534), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n535), .A2(n545), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n536), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n539) );
  NAND2_X1 U609 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U610 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n545), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n543), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n546), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U616 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(KEYINPUT54), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT119), .B(n548), .ZN(n549) );
  NOR2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n573) );
  NAND2_X1 U622 ( .A1(n555), .A2(n573), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT55), .B(n556), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n569) );
  NOR2_X1 U625 ( .A1(n574), .A2(n569), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT122), .B(n559), .Z(n560) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n569), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n564), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n569), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G190GAT), .B(n570), .Z(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT58), .B(n571), .ZN(G1351GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n574), .A2(n584), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  INV_X1 U643 ( .A(n584), .ZN(n588) );
  AND2_X1 U644 ( .A1(n578), .A2(n588), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(KEYINPUT124), .B(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

