

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784;

  OR2_X1 U369 ( .A1(n415), .A2(n412), .ZN(n673) );
  OR2_X1 U370 ( .A1(n648), .A2(G902), .ZN(n514) );
  XNOR2_X1 U371 ( .A(n479), .B(n478), .ZN(n500) );
  XNOR2_X1 U372 ( .A(n455), .B(n468), .ZN(n480) );
  XNOR2_X1 U373 ( .A(G146), .B(G125), .ZN(n467) );
  NOR2_X2 U374 ( .A1(n598), .A2(n747), .ZN(n616) );
  XNOR2_X1 U375 ( .A(G119), .B(G128), .ZN(n516) );
  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n504) );
  AND2_X1 U377 ( .A1(n664), .A2(KEYINPUT81), .ZN(n665) );
  NOR2_X1 U378 ( .A1(n368), .A2(n367), .ZN(n372) );
  INV_X2 U379 ( .A(G953), .ZN(n775) );
  XNOR2_X2 U380 ( .A(n629), .B(n628), .ZN(n634) );
  NOR2_X2 U381 ( .A1(n586), .A2(n575), .ZN(n572) );
  AND2_X2 U382 ( .A1(n365), .A2(n375), .ZN(n374) );
  AND2_X2 U383 ( .A1(n378), .A2(n596), .ZN(n534) );
  NAND2_X1 U384 ( .A1(n417), .A2(n713), .ZN(n414) );
  NAND2_X1 U385 ( .A1(n425), .A2(n424), .ZN(n430) );
  AND2_X1 U386 ( .A1(n426), .A2(n350), .ZN(n425) );
  XNOR2_X1 U387 ( .A(n546), .B(n377), .ZN(n379) );
  XNOR2_X1 U388 ( .A(n438), .B(n503), .ZN(n546) );
  XNOR2_X1 U389 ( .A(n491), .B(n490), .ZN(n672) );
  XNOR2_X1 U390 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U391 ( .A(KEYINPUT20), .B(n489), .ZN(n524) );
  XNOR2_X1 U392 ( .A(n456), .B(KEYINPUT15), .ZN(n626) );
  XNOR2_X2 U393 ( .A(n573), .B(KEYINPUT40), .ZN(n783) );
  AND2_X1 U394 ( .A1(n672), .A2(KEYINPUT68), .ZN(n411) );
  XNOR2_X2 U395 ( .A(n421), .B(n420), .ZN(n782) );
  NOR2_X1 U396 ( .A1(n530), .A2(n596), .ZN(n541) );
  XNOR2_X2 U397 ( .A(n423), .B(n509), .ZN(n756) );
  NAND2_X2 U398 ( .A1(n361), .A2(n407), .ZN(n679) );
  NOR2_X1 U399 ( .A1(n402), .A2(n401), .ZN(n361) );
  XNOR2_X1 U400 ( .A(n581), .B(n529), .ZN(n596) );
  NAND2_X1 U401 ( .A1(n727), .A2(n502), .ZN(n438) );
  AND2_X1 U402 ( .A1(n415), .A2(n411), .ZN(n401) );
  XNOR2_X1 U403 ( .A(n488), .B(KEYINPUT107), .ZN(n574) );
  XNOR2_X1 U404 ( .A(n467), .B(KEYINPUT10), .ZN(n769) );
  NAND2_X1 U405 ( .A1(n356), .A2(n539), .ZN(n355) );
  INV_X1 U406 ( .A(n718), .ZN(n356) );
  NAND2_X1 U407 ( .A1(n440), .A2(n358), .ZN(n538) );
  INV_X1 U408 ( .A(n782), .ZN(n358) );
  XNOR2_X1 U409 ( .A(G113), .B(G101), .ZN(n453) );
  XOR2_X1 U410 ( .A(G110), .B(G137), .Z(n517) );
  XNOR2_X1 U411 ( .A(n387), .B(n388), .ZN(n386) );
  XNOR2_X1 U412 ( .A(n390), .B(n389), .ZN(n388) );
  XNOR2_X1 U413 ( .A(n385), .B(n384), .ZN(n387) );
  XNOR2_X1 U414 ( .A(G143), .B(G104), .ZN(n469) );
  XOR2_X1 U415 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n470) );
  XNOR2_X1 U416 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U417 ( .A(n480), .B(n347), .ZN(n423) );
  XNOR2_X1 U418 ( .A(n772), .B(G146), .ZN(n511) );
  NAND2_X1 U419 ( .A1(n370), .A2(KEYINPUT35), .ZN(n369) );
  NOR2_X1 U420 ( .A1(n678), .A2(KEYINPUT108), .ZN(n428) );
  INV_X1 U421 ( .A(n673), .ZN(n441) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n377) );
  XNOR2_X1 U423 ( .A(n523), .B(n522), .ZN(n713) );
  XNOR2_X1 U424 ( .A(n521), .B(n348), .ZN(n522) );
  XNOR2_X1 U425 ( .A(n400), .B(n399), .ZN(n523) );
  XNOR2_X1 U426 ( .A(G113), .B(KEYINPUT12), .ZN(n384) );
  XNOR2_X1 U427 ( .A(G140), .B(KEYINPUT102), .ZN(n385) );
  XNOR2_X1 U428 ( .A(G122), .B(KEYINPUT11), .ZN(n390) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT90), .ZN(n456) );
  NOR2_X1 U430 ( .A1(KEYINPUT4), .A2(G953), .ZN(n444) );
  NAND2_X1 U431 ( .A1(n443), .A2(G224), .ZN(n442) );
  INV_X1 U432 ( .A(G953), .ZN(n443) );
  XNOR2_X1 U433 ( .A(n355), .B(KEYINPUT67), .ZN(n354) );
  INV_X1 U434 ( .A(KEYINPUT86), .ZN(n360) );
  OR2_X1 U435 ( .A1(G237), .A2(G902), .ZN(n459) );
  NAND2_X1 U436 ( .A1(n410), .A2(n408), .ZN(n402) );
  NAND2_X1 U437 ( .A1(n409), .A2(n531), .ZN(n408) );
  NOR2_X1 U438 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U439 ( .A1(n417), .A2(G902), .ZN(n413) );
  XNOR2_X1 U440 ( .A(n453), .B(n452), .ZN(n422) );
  INV_X1 U441 ( .A(KEYINPUT72), .ZN(n452) );
  XNOR2_X1 U442 ( .A(n500), .B(n499), .ZN(n772) );
  XNOR2_X1 U443 ( .A(KEYINPUT4), .B(G137), .ZN(n498) );
  XNOR2_X1 U444 ( .A(G131), .B(KEYINPUT70), .ZN(n497) );
  XNOR2_X1 U445 ( .A(n437), .B(KEYINPUT69), .ZN(n520) );
  INV_X1 U446 ( .A(G140), .ZN(n437) );
  XNOR2_X1 U447 ( .A(n451), .B(n393), .ZN(n392) );
  INV_X1 U448 ( .A(KEYINPUT73), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n349), .B(n448), .ZN(n449) );
  XNOR2_X1 U450 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n448) );
  XOR2_X1 U451 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n349) );
  NOR2_X1 U452 ( .A1(n433), .A2(n435), .ZN(n431) );
  INV_X1 U453 ( .A(n588), .ZN(n435) );
  AND2_X1 U454 ( .A1(n536), .A2(n352), .ZN(n434) );
  NAND2_X1 U455 ( .A1(n528), .A2(n502), .ZN(n416) );
  XNOR2_X1 U456 ( .A(n518), .B(n515), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n517), .B(n516), .ZN(n518) );
  INV_X1 U458 ( .A(n769), .ZN(n399) );
  INV_X1 U459 ( .A(G134), .ZN(n478) );
  XNOR2_X1 U460 ( .A(n471), .B(n447), .ZN(n472) );
  XNOR2_X1 U461 ( .A(n386), .B(n769), .ZN(n473) );
  XNOR2_X1 U462 ( .A(n520), .B(n436), .ZN(n770) );
  INV_X1 U463 ( .A(KEYINPUT94), .ZN(n436) );
  XOR2_X1 U464 ( .A(G101), .B(G107), .Z(n495) );
  INV_X1 U465 ( .A(KEYINPUT91), .ZN(n450) );
  NAND2_X1 U466 ( .A1(G234), .A2(G237), .ZN(n462) );
  NAND2_X1 U467 ( .A1(n692), .A2(n380), .ZN(n694) );
  NOR2_X1 U468 ( .A1(n662), .A2(KEYINPUT81), .ZN(n668) );
  XOR2_X1 U469 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  XNOR2_X1 U470 ( .A(n655), .B(KEYINPUT59), .ZN(n656) );
  XNOR2_X1 U471 ( .A(n501), .B(n511), .ZN(n727) );
  XNOR2_X1 U472 ( .A(n364), .B(n362), .ZN(n501) );
  XNOR2_X1 U473 ( .A(n757), .B(KEYINPUT73), .ZN(n362) );
  XNOR2_X1 U474 ( .A(n770), .B(n496), .ZN(n364) );
  XNOR2_X1 U475 ( .A(n636), .B(n639), .ZN(n640) );
  XNOR2_X1 U476 ( .A(n585), .B(n383), .ZN(n784) );
  OR2_X1 U477 ( .A1(n604), .A2(n379), .ZN(n647) );
  NAND2_X1 U478 ( .A1(n372), .A2(n376), .ZN(n371) );
  INV_X1 U479 ( .A(G122), .ZN(n468) );
  INV_X1 U480 ( .A(KEYINPUT32), .ZN(n420) );
  AND2_X1 U481 ( .A1(n678), .A2(n441), .ZN(n439) );
  OR2_X1 U482 ( .A1(n618), .A2(n586), .ZN(n587) );
  NOR2_X1 U483 ( .A1(n592), .A2(n591), .ZN(n745) );
  XOR2_X1 U484 ( .A(n713), .B(KEYINPUT122), .Z(n714) );
  INV_X1 U485 ( .A(n379), .ZN(n678) );
  XNOR2_X1 U486 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n347) );
  XOR2_X1 U487 ( .A(n520), .B(KEYINPUT95), .Z(n348) );
  BUF_X1 U488 ( .A(n630), .Z(n663) );
  AND2_X1 U489 ( .A1(n427), .A2(n581), .ZN(n350) );
  INV_X1 U490 ( .A(G902), .ZN(n502) );
  INV_X1 U491 ( .A(n440), .ZN(n739) );
  XOR2_X1 U492 ( .A(n465), .B(KEYINPUT0), .Z(n351) );
  XOR2_X1 U493 ( .A(KEYINPUT78), .B(KEYINPUT34), .Z(n352) );
  XOR2_X1 U494 ( .A(KEYINPUT84), .B(KEYINPUT46), .Z(n353) );
  XNOR2_X1 U495 ( .A(n419), .B(n467), .ZN(n418) );
  NAND2_X1 U496 ( .A1(n445), .A2(n446), .ZN(n419) );
  BUF_X1 U497 ( .A(n719), .Z(n725) );
  NAND2_X1 U498 ( .A1(n434), .A2(n705), .ZN(n432) );
  XNOR2_X2 U499 ( .A(n534), .B(n533), .ZN(n705) );
  NAND2_X1 U500 ( .A1(n406), .A2(n403), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n538), .B(n360), .ZN(n357) );
  NAND2_X1 U502 ( .A1(n357), .A2(n354), .ZN(n359) );
  NAND2_X1 U503 ( .A1(n396), .A2(n441), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n359), .B(KEYINPUT74), .ZN(n559) );
  XNOR2_X1 U505 ( .A(n392), .B(n449), .ZN(n391) );
  NAND2_X1 U506 ( .A1(n442), .A2(KEYINPUT4), .ZN(n446) );
  INV_X1 U507 ( .A(n528), .ZN(n417) );
  NAND2_X1 U508 ( .A1(n444), .A2(G224), .ZN(n445) );
  XNOR2_X2 U509 ( .A(G116), .B(G107), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n395), .B(n756), .ZN(n635) );
  XNOR2_X2 U511 ( .A(n363), .B(n450), .ZN(n757) );
  XNOR2_X2 U512 ( .A(G110), .B(G104), .ZN(n363) );
  NAND2_X1 U513 ( .A1(n366), .A2(KEYINPUT35), .ZN(n365) );
  NAND2_X1 U514 ( .A1(n432), .A2(n431), .ZN(n366) );
  INV_X1 U515 ( .A(n432), .ZN(n367) );
  NAND2_X1 U516 ( .A1(n431), .A2(n373), .ZN(n368) );
  OR2_X1 U517 ( .A1(n705), .A2(n352), .ZN(n376) );
  OR2_X1 U518 ( .A1(n705), .A2(n369), .ZN(n375) );
  INV_X1 U519 ( .A(n352), .ZN(n370) );
  NAND2_X2 U520 ( .A1(n374), .A2(n371), .ZN(n718) );
  INV_X1 U521 ( .A(KEYINPUT35), .ZN(n373) );
  NOR2_X1 U522 ( .A1(n532), .A2(n379), .ZN(n378) );
  XNOR2_X2 U523 ( .A(n514), .B(n513), .ZN(n581) );
  INV_X1 U524 ( .A(n574), .ZN(n380) );
  NAND2_X1 U525 ( .A1(n611), .A2(n381), .ZN(n613) );
  XNOR2_X1 U526 ( .A(n382), .B(n353), .ZN(n381) );
  NAND2_X1 U527 ( .A1(n784), .A2(n783), .ZN(n382) );
  INV_X1 U528 ( .A(KEYINPUT42), .ZN(n383) );
  INV_X1 U529 ( .A(G131), .ZN(n389) );
  XNOR2_X1 U530 ( .A(n394), .B(n391), .ZN(n395) );
  XNOR2_X1 U531 ( .A(n418), .B(n757), .ZN(n394) );
  AND2_X2 U532 ( .A1(n634), .A2(n633), .ZN(n719) );
  XNOR2_X1 U533 ( .A(n430), .B(KEYINPUT65), .ZN(n396) );
  NAND2_X1 U534 ( .A1(n429), .A2(n428), .ZN(n424) );
  XNOR2_X1 U535 ( .A(n560), .B(KEYINPUT45), .ZN(n630) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n655) );
  XNOR2_X2 U537 ( .A(G143), .B(G128), .ZN(n479) );
  INV_X1 U538 ( .A(n397), .ZN(n398) );
  NAND2_X1 U539 ( .A1(n630), .A2(n397), .ZN(n625) );
  AND2_X2 U540 ( .A1(n624), .A2(n623), .ZN(n397) );
  NAND2_X1 U541 ( .A1(n397), .A2(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U542 ( .A1(n397), .A2(n665), .ZN(n666) );
  XNOR2_X1 U543 ( .A(n398), .B(n777), .ZN(n776) );
  NAND2_X1 U544 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U545 ( .A1(n413), .A2(n531), .ZN(n404) );
  INV_X1 U546 ( .A(n414), .ZN(n405) );
  INV_X1 U547 ( .A(n415), .ZN(n406) );
  INV_X1 U548 ( .A(n672), .ZN(n409) );
  NAND2_X1 U549 ( .A1(n412), .A2(n411), .ZN(n410) );
  NOR2_X1 U550 ( .A1(n416), .A2(n713), .ZN(n415) );
  NAND2_X1 U551 ( .A1(n541), .A2(n439), .ZN(n421) );
  XNOR2_X2 U552 ( .A(n422), .B(n454), .ZN(n509) );
  INV_X1 U553 ( .A(n530), .ZN(n429) );
  NAND2_X1 U554 ( .A1(n530), .A2(KEYINPUT108), .ZN(n426) );
  NAND2_X1 U555 ( .A1(n678), .A2(KEYINPUT108), .ZN(n427) );
  NOR2_X1 U556 ( .A1(n536), .A2(n352), .ZN(n433) );
  INV_X1 U557 ( .A(n669), .ZN(n633) );
  AND2_X1 U558 ( .A1(G214), .A2(n504), .ZN(n447) );
  XNOR2_X1 U559 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n515) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n628) );
  XNOR2_X1 U561 ( .A(n477), .B(n476), .ZN(n537) );
  INV_X1 U562 ( .A(n479), .ZN(n451) );
  XOR2_X1 U563 ( .A(KEYINPUT3), .B(G119), .Z(n454) );
  NAND2_X1 U564 ( .A1(n635), .A2(n626), .ZN(n458) );
  AND2_X1 U565 ( .A1(n459), .A2(G210), .ZN(n457) );
  XNOR2_X2 U566 ( .A(n458), .B(n457), .ZN(n569) );
  NAND2_X1 U567 ( .A1(G214), .A2(n459), .ZN(n691) );
  NAND2_X1 U568 ( .A1(n569), .A2(n691), .ZN(n599) );
  INV_X1 U569 ( .A(KEYINPUT19), .ZN(n460) );
  XNOR2_X1 U570 ( .A(n599), .B(n460), .ZN(n590) );
  NOR2_X1 U571 ( .A1(G898), .A2(n775), .ZN(n759) );
  NAND2_X1 U572 ( .A1(n759), .A2(G902), .ZN(n461) );
  NAND2_X1 U573 ( .A1(G952), .A2(n775), .ZN(n562) );
  NAND2_X1 U574 ( .A1(n461), .A2(n562), .ZN(n463) );
  XNOR2_X1 U575 ( .A(n462), .B(KEYINPUT14), .ZN(n701) );
  NAND2_X1 U576 ( .A1(n463), .A2(n701), .ZN(n464) );
  NOR2_X2 U577 ( .A1(n590), .A2(n464), .ZN(n466) );
  INV_X1 U578 ( .A(KEYINPUT66), .ZN(n465) );
  XNOR2_X1 U579 ( .A(n466), .B(n351), .ZN(n535) );
  XNOR2_X1 U580 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U581 ( .A1(G902), .A2(n655), .ZN(n477) );
  XNOR2_X1 U582 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n475) );
  INV_X1 U583 ( .A(G475), .ZN(n474) );
  XNOR2_X1 U584 ( .A(n480), .B(n500), .ZN(n485) );
  XOR2_X1 U585 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n483) );
  NAND2_X1 U586 ( .A1(G234), .A2(n775), .ZN(n481) );
  XOR2_X1 U587 ( .A(KEYINPUT8), .B(n481), .Z(n519) );
  NAND2_X1 U588 ( .A1(G217), .A2(n519), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U590 ( .A(n485), .B(n484), .ZN(n720) );
  NAND2_X1 U591 ( .A1(n720), .A2(n502), .ZN(n487) );
  INV_X1 U592 ( .A(G478), .ZN(n486) );
  XNOR2_X1 U593 ( .A(n487), .B(n486), .ZN(n551) );
  NAND2_X1 U594 ( .A1(n537), .A2(n551), .ZN(n488) );
  NAND2_X1 U595 ( .A1(n626), .A2(G234), .ZN(n489) );
  NAND2_X1 U596 ( .A1(n524), .A2(G221), .ZN(n491) );
  XNOR2_X1 U597 ( .A(KEYINPUT97), .B(KEYINPUT21), .ZN(n490) );
  AND2_X1 U598 ( .A1(n574), .A2(n672), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n535), .A2(n492), .ZN(n493) );
  XNOR2_X2 U600 ( .A(n493), .B(KEYINPUT22), .ZN(n530) );
  NAND2_X1 U601 ( .A1(G227), .A2(n775), .ZN(n494) );
  XNOR2_X1 U602 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U603 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U604 ( .A(KEYINPUT71), .B(G469), .Z(n503) );
  NAND2_X1 U605 ( .A1(n504), .A2(G210), .ZN(n505) );
  XNOR2_X1 U606 ( .A(n505), .B(G116), .ZN(n507) );
  XNOR2_X1 U607 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U609 ( .A(n508), .B(n509), .ZN(n510) );
  XNOR2_X1 U610 ( .A(n511), .B(n510), .ZN(n648) );
  INV_X1 U611 ( .A(KEYINPUT100), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n512), .B(G472), .ZN(n513) );
  NAND2_X1 U613 ( .A1(n519), .A2(G221), .ZN(n521) );
  NAND2_X1 U614 ( .A1(n524), .A2(G217), .ZN(n527) );
  XNOR2_X1 U615 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n525) );
  XOR2_X1 U616 ( .A(n525), .B(KEYINPUT96), .Z(n526) );
  XNOR2_X1 U617 ( .A(KEYINPUT106), .B(KEYINPUT6), .ZN(n529) );
  INV_X1 U618 ( .A(KEYINPUT68), .ZN(n531) );
  INV_X1 U619 ( .A(n679), .ZN(n532) );
  XNOR2_X1 U620 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n533) );
  BUF_X1 U621 ( .A(n535), .Z(n536) );
  NOR2_X1 U622 ( .A1(n537), .A2(n551), .ZN(n588) );
  NOR2_X1 U623 ( .A1(n538), .A2(n718), .ZN(n540) );
  INV_X1 U624 ( .A(KEYINPUT44), .ZN(n539) );
  NOR2_X1 U625 ( .A1(n540), .A2(n539), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n541), .B(KEYINPUT85), .ZN(n543) );
  NAND2_X1 U627 ( .A1(n673), .A2(n379), .ZN(n542) );
  OR2_X1 U628 ( .A1(n543), .A2(n542), .ZN(n732) );
  INV_X1 U629 ( .A(n536), .ZN(n547) );
  NOR2_X1 U630 ( .A1(n379), .A2(n581), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n679), .A2(n544), .ZN(n684) );
  NOR2_X1 U632 ( .A1(n547), .A2(n684), .ZN(n545) );
  XNOR2_X1 U633 ( .A(n545), .B(KEYINPUT31), .ZN(n749) );
  NAND2_X1 U634 ( .A1(n546), .A2(n679), .ZN(n565) );
  NOR2_X1 U635 ( .A1(n565), .A2(n547), .ZN(n548) );
  XNOR2_X1 U636 ( .A(KEYINPUT98), .B(n548), .ZN(n549) );
  NAND2_X1 U637 ( .A1(n549), .A2(n581), .ZN(n736) );
  NAND2_X1 U638 ( .A1(n749), .A2(n736), .ZN(n554) );
  INV_X1 U639 ( .A(KEYINPUT105), .ZN(n550) );
  XNOR2_X1 U640 ( .A(n537), .B(n550), .ZN(n553) );
  INV_X1 U641 ( .A(n551), .ZN(n552) );
  NAND2_X1 U642 ( .A1(n553), .A2(n552), .ZN(n750) );
  OR2_X1 U643 ( .A1(n553), .A2(n552), .ZN(n747) );
  NAND2_X1 U644 ( .A1(n750), .A2(n747), .ZN(n690) );
  NAND2_X1 U645 ( .A1(n554), .A2(n690), .ZN(n555) );
  NAND2_X1 U646 ( .A1(n732), .A2(n555), .ZN(n556) );
  NOR2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U648 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U649 ( .A(n747), .ZN(n744) );
  NOR2_X1 U650 ( .A1(G900), .A2(n775), .ZN(n561) );
  NAND2_X1 U651 ( .A1(n561), .A2(G902), .ZN(n563) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U653 ( .A1(n564), .A2(n701), .ZN(n578) );
  NOR2_X1 U654 ( .A1(n578), .A2(n565), .ZN(n568) );
  INV_X1 U655 ( .A(n691), .ZN(n614) );
  NOR2_X1 U656 ( .A1(n581), .A2(n614), .ZN(n566) );
  XNOR2_X1 U657 ( .A(n566), .B(KEYINPUT30), .ZN(n567) );
  NAND2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n586) );
  BUF_X1 U659 ( .A(n569), .Z(n570) );
  XOR2_X1 U660 ( .A(KEYINPUT38), .B(n570), .Z(n693) );
  INV_X1 U661 ( .A(n693), .ZN(n575) );
  INV_X1 U662 ( .A(KEYINPUT39), .ZN(n571) );
  XNOR2_X1 U663 ( .A(n572), .B(n571), .ZN(n622) );
  NAND2_X1 U664 ( .A1(n744), .A2(n622), .ZN(n573) );
  NAND2_X1 U665 ( .A1(n574), .A2(n691), .ZN(n696) );
  NOR2_X1 U666 ( .A1(n575), .A2(n696), .ZN(n577) );
  XOR2_X1 U667 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n576) );
  XNOR2_X1 U668 ( .A(n577), .B(n576), .ZN(n688) );
  INV_X1 U669 ( .A(n578), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n672), .A2(n579), .ZN(n580) );
  NOR2_X1 U671 ( .A1(n673), .A2(n580), .ZN(n597) );
  INV_X1 U672 ( .A(n581), .ZN(n675) );
  NAND2_X1 U673 ( .A1(n597), .A2(n675), .ZN(n583) );
  XOR2_X1 U674 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n582) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n584), .A2(n546), .ZN(n592) );
  NOR2_X1 U677 ( .A1(n688), .A2(n592), .ZN(n585) );
  INV_X1 U678 ( .A(n570), .ZN(n618) );
  XNOR2_X1 U679 ( .A(KEYINPUT109), .B(n587), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n743) );
  BUF_X1 U681 ( .A(n590), .Z(n591) );
  NAND2_X1 U682 ( .A1(n690), .A2(n745), .ZN(n593) );
  NAND2_X1 U683 ( .A1(n593), .A2(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U684 ( .A1(n743), .A2(n594), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n595), .B(KEYINPUT80), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT112), .ZN(n602) );
  BUF_X1 U688 ( .A(n599), .Z(n600) );
  INV_X1 U689 ( .A(n600), .ZN(n601) );
  NAND2_X1 U690 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT36), .ZN(n604) );
  INV_X1 U692 ( .A(n690), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n605), .A2(KEYINPUT47), .ZN(n606) );
  XNOR2_X1 U694 ( .A(n606), .B(KEYINPUT76), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n745), .A2(n607), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n647), .A2(n608), .ZN(n609) );
  NOR2_X1 U697 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U698 ( .A(KEYINPUT48), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n613), .B(n612), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n678), .A2(n614), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U702 ( .A(n617), .B(KEYINPUT43), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n754) );
  NAND2_X1 U704 ( .A1(n620), .A2(n754), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT83), .ZN(n624) );
  INV_X1 U706 ( .A(n750), .ZN(n740) );
  AND2_X1 U707 ( .A1(n622), .A2(n740), .ZN(n752) );
  INV_X1 U708 ( .A(n752), .ZN(n623) );
  INV_X1 U709 ( .A(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U710 ( .A1(n625), .A2(n664), .ZN(n661) );
  INV_X1 U711 ( .A(n626), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n661), .A2(n627), .ZN(n629) );
  INV_X1 U713 ( .A(n663), .ZN(n632) );
  NOR2_X2 U714 ( .A1(n632), .A2(n631), .ZN(n669) );
  NAND2_X1 U715 ( .A1(n719), .A2(G210), .ZN(n641) );
  BUF_X1 U716 ( .A(n635), .Z(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n638) );
  XNOR2_X1 U718 ( .A(KEYINPUT88), .B(KEYINPUT79), .ZN(n637) );
  XOR2_X1 U719 ( .A(n638), .B(n637), .Z(n639) );
  XNOR2_X1 U720 ( .A(n641), .B(n640), .ZN(n643) );
  INV_X1 U721 ( .A(G952), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n642), .A2(G953), .ZN(n723) );
  NAND2_X1 U723 ( .A1(n643), .A2(n723), .ZN(n645) );
  INV_X1 U724 ( .A(KEYINPUT56), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n645), .B(n644), .ZN(G51) );
  XOR2_X1 U726 ( .A(G125), .B(KEYINPUT37), .Z(n646) );
  XNOR2_X1 U727 ( .A(n647), .B(n646), .ZN(G27) );
  NAND2_X1 U728 ( .A1(n719), .A2(G472), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n651), .A2(n723), .ZN(n654) );
  XNOR2_X1 U731 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(KEYINPUT87), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n654), .B(n653), .ZN(G57) );
  NAND2_X1 U734 ( .A1(n719), .A2(G475), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n658), .A2(n723), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT120), .B(KEYINPUT60), .Z(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(G60) );
  INV_X1 U739 ( .A(n661), .ZN(n662) );
  NOR2_X1 U740 ( .A1(n663), .A2(n666), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT82), .B(n671), .Z(n710) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U745 ( .A(KEYINPUT49), .B(n674), .Z(n676) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT117), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n680), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n683), .B(KEYINPUT118), .ZN(n686) );
  INV_X1 U752 ( .A(n684), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n687), .ZN(n689) );
  INV_X1 U755 ( .A(n688), .ZN(n704) );
  NAND2_X1 U756 ( .A1(n689), .A2(n704), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n705), .A2(n697), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U762 ( .A(KEYINPUT52), .B(n700), .Z(n703) );
  NAND2_X1 U763 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n708) );
  NAND2_X1 U765 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U766 ( .A1(n706), .A2(n775), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U768 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U769 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n711) );
  XNOR2_X1 U770 ( .A(n712), .B(n711), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n719), .A2(G217), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n716), .A2(n723), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n717), .B(KEYINPUT123), .ZN(G66) );
  XNOR2_X1 U775 ( .A(n718), .B(n468), .ZN(G24) );
  NAND2_X1 U776 ( .A1(n725), .A2(G478), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n720), .B(KEYINPUT121), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(n724) );
  INV_X1 U779 ( .A(n723), .ZN(n730) );
  NOR2_X1 U780 ( .A1(n724), .A2(n730), .ZN(G63) );
  NAND2_X1 U781 ( .A1(n725), .A2(G469), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n731) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(G54) );
  XNOR2_X1 U786 ( .A(G101), .B(n732), .ZN(G3) );
  NOR2_X1 U787 ( .A1(n736), .A2(n747), .ZN(n733) );
  XOR2_X1 U788 ( .A(G104), .B(n733), .Z(G6) );
  XOR2_X1 U789 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n735) );
  XNOR2_X1 U790 ( .A(G107), .B(KEYINPUT27), .ZN(n734) );
  XNOR2_X1 U791 ( .A(n735), .B(n734), .ZN(n738) );
  NOR2_X1 U792 ( .A1(n736), .A2(n750), .ZN(n737) );
  XOR2_X1 U793 ( .A(n738), .B(n737), .Z(G9) );
  XOR2_X1 U794 ( .A(n739), .B(G110), .Z(G12) );
  XOR2_X1 U795 ( .A(G128), .B(KEYINPUT29), .Z(n742) );
  NAND2_X1 U796 ( .A1(n745), .A2(n740), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n742), .B(n741), .ZN(G30) );
  XNOR2_X1 U798 ( .A(n743), .B(G143), .ZN(G45) );
  NAND2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n746), .B(G146), .ZN(G48) );
  NOR2_X1 U801 ( .A1(n747), .A2(n749), .ZN(n748) );
  XOR2_X1 U802 ( .A(G113), .B(n748), .Z(G15) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U804 ( .A(G116), .B(n751), .Z(G18) );
  XNOR2_X1 U805 ( .A(G134), .B(n752), .ZN(n753) );
  XNOR2_X1 U806 ( .A(n753), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U807 ( .A(G140), .B(KEYINPUT116), .ZN(n755) );
  XNOR2_X1 U808 ( .A(n755), .B(n754), .ZN(G42) );
  XNOR2_X1 U809 ( .A(n756), .B(n757), .ZN(n758) );
  NOR2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(KEYINPUT126), .B(n760), .ZN(n768) );
  NAND2_X1 U812 ( .A1(G224), .A2(G953), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n761), .B(KEYINPUT61), .ZN(n762) );
  XNOR2_X1 U814 ( .A(KEYINPUT124), .B(n762), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n763), .A2(G898), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n663), .A2(n775), .ZN(n764) );
  XOR2_X1 U817 ( .A(KEYINPUT125), .B(n764), .Z(n765) );
  NAND2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(G69) );
  XOR2_X1 U820 ( .A(KEYINPUT127), .B(n769), .Z(n771) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n774) );
  INV_X1 U822 ( .A(n772), .ZN(n773) );
  XNOR2_X1 U823 ( .A(n774), .B(n773), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n776), .A2(n775), .ZN(n781) );
  XNOR2_X1 U825 ( .A(G227), .B(n777), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(G900), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n779), .A2(G953), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n781), .A2(n780), .ZN(G72) );
  XOR2_X1 U829 ( .A(G119), .B(n782), .Z(G21) );
  XNOR2_X1 U830 ( .A(G131), .B(n783), .ZN(G33) );
  XNOR2_X1 U831 ( .A(G137), .B(n784), .ZN(G39) );
endmodule

