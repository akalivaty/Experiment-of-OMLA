

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U558 ( .A1(G8), .A2(n669), .ZN(n703) );
  XNOR2_X1 U559 ( .A(G2104), .B(KEYINPUT65), .ZN(n582) );
  AND2_X1 U560 ( .A1(n593), .A2(n592), .ZN(G164) );
  NOR2_X2 U561 ( .A1(G164), .A2(G1384), .ZN(n711) );
  BUF_X1 U562 ( .A(n995), .Z(n524) );
  BUF_X1 U563 ( .A(n995), .Z(n525) );
  NOR2_X1 U564 ( .A1(G2105), .A2(n582), .ZN(n995) );
  AND2_X1 U565 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U566 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X2 U567 ( .A1(n587), .A2(n586), .ZN(G160) );
  INV_X1 U568 ( .A(KEYINPUT28), .ZN(n657) );
  XNOR2_X1 U569 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n599) );
  NOR2_X1 U570 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U571 ( .A1(n703), .A2(n691), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n649), .B(KEYINPUT94), .ZN(n650) );
  XNOR2_X1 U573 ( .A(n651), .B(n650), .ZN(n653) );
  XNOR2_X1 U574 ( .A(n600), .B(n599), .ZN(n601) );
  NOR2_X2 U575 ( .A1(n710), .A2(n594), .ZN(n616) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n567) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U578 ( .A1(G86), .A2(n791), .ZN(n529) );
  NOR2_X1 U579 ( .A1(G651), .A2(n567), .ZN(n527) );
  XNOR2_X2 U580 ( .A(KEYINPUT64), .B(n527), .ZN(n796) );
  NAND2_X1 U581 ( .A1(G48), .A2(n796), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n532) );
  INV_X1 U583 ( .A(G651), .ZN(n533) );
  NOR2_X1 U584 ( .A1(n567), .A2(n533), .ZN(n792) );
  NAND2_X1 U585 ( .A1(n792), .A2(G73), .ZN(n530) );
  XOR2_X1 U586 ( .A(KEYINPUT2), .B(n530), .Z(n531) );
  NOR2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X2 U589 ( .A(KEYINPUT1), .B(n534), .Z(n795) );
  NAND2_X1 U590 ( .A1(n795), .A2(G61), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(G305) );
  NAND2_X1 U592 ( .A1(n791), .A2(G89), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n537), .B(KEYINPUT4), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G76), .A2(n792), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT5), .ZN(n547) );
  XNOR2_X1 U597 ( .A(KEYINPUT73), .B(KEYINPUT6), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G51), .A2(n796), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT72), .ZN(n543) );
  NAND2_X1 U600 ( .A1(G63), .A2(n795), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U604 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  NAND2_X1 U605 ( .A1(n795), .A2(G64), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G52), .A2(n796), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U608 ( .A1(G90), .A2(n791), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G77), .A2(n792), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U613 ( .A(G171), .ZN(G301) );
  XOR2_X1 U614 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U615 ( .A1(n795), .A2(G62), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G50), .A2(n796), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G88), .A2(n791), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G75), .A2(n792), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U622 ( .A(n562), .B(KEYINPUT77), .Z(G166) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(G651), .A2(G74), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G49), .A2(n796), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U627 ( .A(KEYINPUT76), .B(n565), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n795), .A2(n566), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n567), .A2(G87), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(G288) );
  AND2_X1 U631 ( .A1(G47), .A2(n796), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G85), .A2(n791), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G72), .A2(n792), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n795), .A2(G60), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(G290) );
  XNOR2_X1 U638 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n577) );
  NOR2_X1 U639 ( .A1(G2105), .A2(G2104), .ZN(n576) );
  XNOR2_X2 U640 ( .A(n577), .B(n576), .ZN(n997) );
  NAND2_X1 U641 ( .A1(G137), .A2(n997), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT68), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G101), .A2(n524), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT23), .B(n579), .Z(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n587) );
  AND2_X1 U646 ( .A1(G2105), .A2(G2104), .ZN(n991) );
  NAND2_X1 U647 ( .A1(G113), .A2(n991), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n582), .A2(G2105), .ZN(n583) );
  XOR2_X2 U649 ( .A(KEYINPUT66), .B(n583), .Z(n992) );
  NAND2_X1 U650 ( .A1(G125), .A2(n992), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n710) );
  NAND2_X1 U653 ( .A1(G102), .A2(n525), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G114), .A2(n991), .ZN(n588) );
  AND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n997), .A2(G138), .ZN(n590) );
  AND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n992), .A2(G126), .ZN(n592) );
  INV_X1 U659 ( .A(n711), .ZN(n594) );
  INV_X1 U660 ( .A(n616), .ZN(n669) );
  NOR2_X1 U661 ( .A1(G1981), .A2(G305), .ZN(n595) );
  XOR2_X1 U662 ( .A(n595), .B(KEYINPUT24), .Z(n596) );
  XNOR2_X1 U663 ( .A(KEYINPUT92), .B(n596), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n703), .A2(n597), .ZN(n708) );
  NOR2_X1 U665 ( .A1(G1966), .A2(n703), .ZN(n679) );
  NOR2_X1 U666 ( .A1(G2084), .A2(n669), .ZN(n681) );
  NOR2_X1 U667 ( .A1(n679), .A2(n681), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G8), .A2(n598), .ZN(n600) );
  NOR2_X1 U669 ( .A1(G168), .A2(n601), .ZN(n605) );
  NAND2_X1 U670 ( .A1(G1961), .A2(n669), .ZN(n603) );
  BUF_X2 U671 ( .A(n616), .Z(n648) );
  XOR2_X1 U672 ( .A(G2078), .B(KEYINPUT25), .Z(n885) );
  NAND2_X1 U673 ( .A1(n648), .A2(n885), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n662) );
  AND2_X1 U675 ( .A1(G301), .A2(n662), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT31), .ZN(n666) );
  NAND2_X1 U678 ( .A1(G56), .A2(n795), .ZN(n607) );
  XOR2_X1 U679 ( .A(KEYINPUT14), .B(n607), .Z(n613) );
  NAND2_X1 U680 ( .A1(n791), .A2(G81), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G68), .A2(n792), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT13), .B(n611), .Z(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G43), .A2(n796), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n1013) );
  NAND2_X1 U688 ( .A1(G1996), .A2(n616), .ZN(n617) );
  XNOR2_X1 U689 ( .A(KEYINPUT26), .B(n617), .ZN(n619) );
  INV_X1 U690 ( .A(G1341), .ZN(n1025) );
  NOR2_X1 U691 ( .A1(n648), .A2(n1025), .ZN(n618) );
  NAND2_X1 U692 ( .A1(KEYINPUT26), .A2(n618), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n619), .A2(n622), .ZN(n621) );
  INV_X1 U694 ( .A(KEYINPUT95), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n622), .A2(KEYINPUT95), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n1013), .A2(n625), .ZN(n637) );
  NAND2_X1 U699 ( .A1(G92), .A2(n791), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G79), .A2(n792), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n795), .A2(G66), .ZN(n629) );
  NAND2_X1 U703 ( .A1(G54), .A2(n796), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U706 ( .A(KEYINPUT15), .B(n632), .Z(n633) );
  XOR2_X2 U707 ( .A(KEYINPUT71), .B(n633), .Z(n1016) );
  INV_X1 U708 ( .A(n1016), .ZN(n639) );
  NAND2_X1 U709 ( .A1(G1348), .A2(n669), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G2067), .A2(n648), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n795), .A2(G65), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G53), .A2(n796), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G91), .A2(n791), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G78), .A2(n792), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n774) );
  NAND2_X1 U722 ( .A1(G2072), .A2(n648), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n649) );
  AND2_X1 U724 ( .A1(G1956), .A2(n669), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n774), .A2(n656), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n774), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT29), .ZN(n664) );
  NOR2_X1 U732 ( .A1(G301), .A2(n662), .ZN(n663) );
  NOR2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n680) );
  INV_X1 U735 ( .A(n680), .ZN(n668) );
  AND2_X1 U736 ( .A1(G286), .A2(G8), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n677) );
  INV_X1 U738 ( .A(G8), .ZN(n675) );
  NOR2_X1 U739 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U740 ( .A(n670), .B(KEYINPUT98), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n703), .A2(G1971), .ZN(n671) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(G303), .ZN(n674) );
  OR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT32), .ZN(n686) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n683) );
  NAND2_X1 U747 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U749 ( .A(n684), .B(KEYINPUT97), .Z(n685) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n702) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n695) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n695), .A2(n687), .ZN(n911) );
  XOR2_X1 U754 ( .A(n911), .B(KEYINPUT99), .Z(n689) );
  INV_X1 U755 ( .A(KEYINPUT33), .ZN(n688) );
  AND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n702), .A2(n690), .ZN(n693) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n910) );
  INV_X1 U759 ( .A(n910), .ZN(n691) );
  OR2_X1 U760 ( .A1(KEYINPUT33), .A2(n526), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n695), .A2(KEYINPUT33), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n703), .A2(n696), .ZN(n697) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U766 ( .A(G1981), .B(G305), .Z(n920) );
  NAND2_X1 U767 ( .A1(n699), .A2(n920), .ZN(n706) );
  NOR2_X1 U768 ( .A1(G2090), .A2(G303), .ZN(n700) );
  NAND2_X1 U769 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n709), .B(KEYINPUT101), .ZN(n748) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n761) );
  XNOR2_X1 U775 ( .A(G1986), .B(G290), .ZN(n906) );
  NAND2_X1 U776 ( .A1(n761), .A2(n906), .ZN(n746) );
  NAND2_X1 U777 ( .A1(G129), .A2(n992), .ZN(n718) );
  NAND2_X1 U778 ( .A1(G141), .A2(n997), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G117), .A2(n991), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n525), .A2(G105), .ZN(n714) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n714), .Z(n715) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U785 ( .A(KEYINPUT89), .B(n719), .Z(n987) );
  NAND2_X1 U786 ( .A1(G1996), .A2(n987), .ZN(n720) );
  XOR2_X1 U787 ( .A(KEYINPUT90), .B(n720), .Z(n728) );
  NAND2_X1 U788 ( .A1(G131), .A2(n997), .ZN(n722) );
  NAND2_X1 U789 ( .A1(G95), .A2(n524), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U791 ( .A1(G107), .A2(n991), .ZN(n724) );
  NAND2_X1 U792 ( .A1(G119), .A2(n992), .ZN(n723) );
  NAND2_X1 U793 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n990) );
  AND2_X1 U795 ( .A1(n990), .A2(G1991), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n865) );
  INV_X1 U797 ( .A(n761), .ZN(n729) );
  NOR2_X1 U798 ( .A1(n865), .A2(n729), .ZN(n753) );
  XOR2_X1 U799 ( .A(KEYINPUT91), .B(n753), .Z(n744) );
  NAND2_X1 U800 ( .A1(G116), .A2(n991), .ZN(n731) );
  NAND2_X1 U801 ( .A1(G128), .A2(n992), .ZN(n730) );
  NAND2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U803 ( .A(KEYINPUT35), .B(n732), .Z(n740) );
  NAND2_X1 U804 ( .A1(n525), .A2(G104), .ZN(n733) );
  XNOR2_X1 U805 ( .A(KEYINPUT85), .B(n733), .ZN(n736) );
  NAND2_X1 U806 ( .A1(n997), .A2(G140), .ZN(n734) );
  XOR2_X1 U807 ( .A(n734), .B(KEYINPUT86), .Z(n735) );
  NOR2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U809 ( .A(KEYINPUT87), .B(n737), .Z(n738) );
  XOR2_X1 U810 ( .A(KEYINPUT34), .B(n738), .Z(n739) );
  NOR2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U812 ( .A(KEYINPUT36), .B(n741), .ZN(n1006) );
  XNOR2_X1 U813 ( .A(G2067), .B(KEYINPUT37), .ZN(n750) );
  NOR2_X1 U814 ( .A1(n1006), .A2(n750), .ZN(n868) );
  NAND2_X1 U815 ( .A1(n868), .A2(n761), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT88), .ZN(n758) );
  INV_X1 U817 ( .A(n758), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT102), .ZN(n764) );
  NAND2_X1 U822 ( .A1(n1006), .A2(n750), .ZN(n873) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n987), .ZN(n861) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n751) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n990), .ZN(n869) );
  NOR2_X1 U826 ( .A1(n751), .A2(n869), .ZN(n752) );
  NOR2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U828 ( .A1(n861), .A2(n754), .ZN(n756) );
  XOR2_X1 U829 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n755) );
  XNOR2_X1 U830 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n873), .A2(n759), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U834 ( .A(n762), .B(KEYINPUT104), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G120), .ZN(G236) );
  INV_X1 U839 ( .A(G69), .ZN(G235) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  XOR2_X1 U843 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n769) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n768) );
  XOR2_X1 U845 ( .A(n769), .B(n768), .Z(n836) );
  INV_X1 U846 ( .A(n836), .ZN(G223) );
  INV_X1 U847 ( .A(G567), .ZN(n831) );
  NOR2_X1 U848 ( .A1(n831), .A2(G223), .ZN(n770) );
  XNOR2_X1 U849 ( .A(n770), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n802) );
  OR2_X1 U851 ( .A1(n1013), .A2(n802), .ZN(G153) );
  NAND2_X1 U852 ( .A1(G301), .A2(G868), .ZN(n771) );
  XNOR2_X1 U853 ( .A(n771), .B(KEYINPUT70), .ZN(n773) );
  OR2_X1 U854 ( .A1(G868), .A2(n1016), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n773), .A2(n772), .ZN(G284) );
  INV_X1 U856 ( .A(n774), .ZN(G299) );
  XOR2_X1 U857 ( .A(KEYINPUT74), .B(G868), .Z(n775) );
  NOR2_X1 U858 ( .A1(G286), .A2(n775), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n802), .A2(G559), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n778), .A2(n1016), .ZN(n779) );
  XNOR2_X1 U863 ( .A(n779), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U864 ( .A1(G868), .A2(n1013), .ZN(n782) );
  NAND2_X1 U865 ( .A1(n1016), .A2(G868), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U868 ( .A1(G135), .A2(n997), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G111), .A2(n991), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n992), .A2(G123), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(KEYINPUT18), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n524), .A2(G99), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n985) );
  XNOR2_X1 U876 ( .A(n985), .B(G2096), .ZN(n790) );
  INV_X1 U877 ( .A(G2100), .ZN(n963) );
  NAND2_X1 U878 ( .A1(n790), .A2(n963), .ZN(G156) );
  NAND2_X1 U879 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n800) );
  NAND2_X1 U882 ( .A1(n795), .A2(G67), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G55), .A2(n796), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n815) );
  NAND2_X1 U886 ( .A1(G559), .A2(n1016), .ZN(n801) );
  XOR2_X1 U887 ( .A(n1013), .B(n801), .Z(n813) );
  NAND2_X1 U888 ( .A1(n802), .A2(n813), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n803), .B(KEYINPUT75), .ZN(n804) );
  XNOR2_X1 U890 ( .A(n815), .B(n804), .ZN(G145) );
  XOR2_X1 U891 ( .A(G303), .B(G305), .Z(n805) );
  XNOR2_X1 U892 ( .A(n805), .B(G288), .ZN(n809) );
  XNOR2_X1 U893 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G290), .B(KEYINPUT19), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n808) );
  XOR2_X1 U896 ( .A(n809), .B(n808), .Z(n811) );
  XOR2_X1 U897 ( .A(G299), .B(n815), .Z(n810) );
  XNOR2_X1 U898 ( .A(n811), .B(n810), .ZN(n1015) );
  XOR2_X1 U899 ( .A(n1015), .B(KEYINPUT80), .Z(n812) );
  XNOR2_X1 U900 ( .A(n813), .B(n812), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n814), .A2(G868), .ZN(n817) );
  OR2_X1 U902 ( .A1(G868), .A2(n815), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U904 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U905 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U906 ( .A1(G2090), .A2(n819), .ZN(n821) );
  XOR2_X1 U907 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G2072), .ZN(n823) );
  XNOR2_X1 U910 ( .A(n823), .B(KEYINPUT82), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n824) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n824), .Z(n825) );
  NOR2_X1 U914 ( .A1(G218), .A2(n825), .ZN(n826) );
  NAND2_X1 U915 ( .A1(G96), .A2(n826), .ZN(n961) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n961), .ZN(n827) );
  XNOR2_X1 U917 ( .A(n827), .B(KEYINPUT83), .ZN(n833) );
  NOR2_X1 U918 ( .A1(G235), .A2(G236), .ZN(n828) );
  XNOR2_X1 U919 ( .A(KEYINPUT84), .B(n828), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n829), .A2(G108), .ZN(n830) );
  NOR2_X1 U921 ( .A1(G237), .A2(n830), .ZN(n960) );
  NOR2_X1 U922 ( .A1(n831), .A2(n960), .ZN(n832) );
  NOR2_X1 U923 ( .A1(n833), .A2(n832), .ZN(G319) );
  INV_X1 U924 ( .A(G319), .ZN(n835) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n834) );
  NOR2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n841) );
  NAND2_X1 U927 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n836), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(n837), .Z(n838) );
  NAND2_X1 U931 ( .A1(n838), .A2(G661), .ZN(n839) );
  XOR2_X1 U932 ( .A(KEYINPUT109), .B(n839), .Z(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n841), .A2(n840), .ZN(G188) );
  XOR2_X1 U935 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  NAND2_X1 U937 ( .A1(G136), .A2(n997), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G112), .A2(n991), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n848) );
  NAND2_X1 U940 ( .A1(n992), .A2(G124), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n525), .A2(G100), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U944 ( .A1(n848), .A2(n847), .ZN(G162) );
  NAND2_X1 U945 ( .A1(G139), .A2(n997), .ZN(n850) );
  NAND2_X1 U946 ( .A1(G103), .A2(n524), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n856) );
  NAND2_X1 U948 ( .A1(G127), .A2(n992), .ZN(n851) );
  XOR2_X1 U949 ( .A(KEYINPUT113), .B(n851), .Z(n853) );
  NAND2_X1 U950 ( .A1(n991), .A2(G115), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT47), .B(n854), .Z(n855) );
  NOR2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n1010) );
  XOR2_X1 U954 ( .A(G2072), .B(n1010), .Z(n858) );
  XOR2_X1 U955 ( .A(G164), .B(G2078), .Z(n857) );
  NOR2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U957 ( .A(KEYINPUT50), .B(n859), .ZN(n864) );
  XOR2_X1 U958 ( .A(G2090), .B(G162), .Z(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT51), .B(n862), .Z(n863) );
  NAND2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n876) );
  XNOR2_X1 U962 ( .A(G160), .B(G2084), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n871) );
  NOR2_X1 U965 ( .A1(n869), .A2(n985), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U967 ( .A(KEYINPUT117), .B(n872), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U969 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U970 ( .A(KEYINPUT52), .B(n877), .ZN(n879) );
  INV_X1 U971 ( .A(KEYINPUT55), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  NAND2_X1 U973 ( .A1(n880), .A2(G29), .ZN(n958) );
  XOR2_X1 U974 ( .A(G34), .B(KEYINPUT120), .Z(n882) );
  XNOR2_X1 U975 ( .A(G2084), .B(KEYINPUT54), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n882), .B(n881), .ZN(n899) );
  XNOR2_X1 U977 ( .A(G2090), .B(G35), .ZN(n897) );
  XNOR2_X1 U978 ( .A(G2067), .B(G26), .ZN(n884) );
  XNOR2_X1 U979 ( .A(G32), .B(G1996), .ZN(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n889) );
  XNOR2_X1 U981 ( .A(n885), .B(G27), .ZN(n887) );
  XNOR2_X1 U982 ( .A(G33), .B(G2072), .ZN(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U985 ( .A(KEYINPUT119), .B(n890), .ZN(n891) );
  NAND2_X1 U986 ( .A1(n891), .A2(G28), .ZN(n894) );
  XNOR2_X1 U987 ( .A(G25), .B(G1991), .ZN(n892) );
  XNOR2_X1 U988 ( .A(KEYINPUT118), .B(n892), .ZN(n893) );
  NOR2_X1 U989 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT53), .B(n895), .ZN(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U993 ( .A(KEYINPUT55), .B(n900), .Z(n902) );
  INV_X1 U994 ( .A(G29), .ZN(n901) );
  NAND2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G11), .A2(n903), .ZN(n956) );
  INV_X1 U997 ( .A(G16), .ZN(n952) );
  XOR2_X1 U998 ( .A(n952), .B(KEYINPUT56), .Z(n928) );
  XNOR2_X1 U999 ( .A(G1961), .B(KEYINPUT122), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n904), .B(G171), .Z(n905) );
  NOR2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n926) );
  XOR2_X1 U1002 ( .A(n1025), .B(KEYINPUT124), .Z(n907) );
  XNOR2_X1 U1003 ( .A(n907), .B(n1013), .ZN(n909) );
  XOR2_X1 U1004 ( .A(G1348), .B(n1016), .Z(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n918) );
  NAND2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G299), .B(G1956), .Z(n913) );
  NAND2_X1 U1008 ( .A1(G1971), .A2(G303), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT123), .B(n916), .Z(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n924) );
  XOR2_X1 U1013 ( .A(G1966), .B(G168), .Z(n919) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(n919), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1016 ( .A(KEYINPUT57), .B(n922), .Z(n923) );
  NOR2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(n928), .A2(n927), .ZN(n954) );
  XOR2_X1 U1020 ( .A(G1976), .B(G23), .Z(n932) );
  XNOR2_X1 U1021 ( .A(G1986), .B(G24), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(G1971), .B(G22), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1025 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(n934), .B(n933), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(G1961), .B(G5), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n948) );
  XOR2_X1 U1031 ( .A(G19), .B(G1341), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G1956), .B(G20), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G6), .B(G1981), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1036 ( .A(KEYINPUT59), .B(G1348), .Z(n943) );
  XNOR2_X1 U1037 ( .A(G4), .B(n943), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1039 ( .A(n946), .B(KEYINPUT60), .Z(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n949), .Z(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT126), .B(n950), .Z(n951) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1046 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1047 ( .A(KEYINPUT62), .B(n959), .Z(G311) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1049 ( .A(G96), .ZN(G221) );
  INV_X1 U1050 ( .A(n960), .ZN(n962) );
  NOR2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(G325) );
  INV_X1 U1052 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1053 ( .A(n963), .B(G2096), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(G2090), .B(KEYINPUT43), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1056 ( .A(n966), .B(KEYINPUT110), .Z(n968) );
  XNOR2_X1 U1057 ( .A(G2072), .B(G2678), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n972) );
  XOR2_X1 U1059 ( .A(KEYINPUT42), .B(G2084), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G2067), .B(G2078), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n972), .B(n971), .ZN(G227) );
  XOR2_X1 U1063 ( .A(G1971), .B(G1961), .Z(n974) );
  XNOR2_X1 U1064 ( .A(G1996), .B(G1966), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n978) );
  XOR2_X1 U1066 ( .A(KEYINPUT111), .B(G2474), .Z(n976) );
  XNOR2_X1 U1067 ( .A(G1991), .B(G1986), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(n978), .B(n977), .Z(n980) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G1976), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n980), .B(n979), .ZN(n982) );
  XOR2_X1 U1072 ( .A(G1981), .B(KEYINPUT41), .Z(n981) );
  XNOR2_X1 U1073 ( .A(n982), .B(n981), .ZN(G229) );
  XOR2_X1 U1074 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G164), .B(KEYINPUT114), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n984), .B(n983), .ZN(n989) );
  XOR2_X1 U1077 ( .A(G160), .B(n985), .Z(n986) );
  XNOR2_X1 U1078 ( .A(n987), .B(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n989), .B(n988), .ZN(n1008) );
  XOR2_X1 U1080 ( .A(n990), .B(G162), .Z(n1004) );
  NAND2_X1 U1081 ( .A1(G118), .A2(n991), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n992), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n1002) );
  NAND2_X1 U1084 ( .A1(n525), .A2(G106), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(n996), .B(KEYINPUT112), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(G142), .A2(n997), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT45), .B(n1000), .Z(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1004), .B(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(n1008), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1093 ( .A(n1010), .B(n1009), .Z(n1011) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1011), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT115), .B(n1012), .Z(G395) );
  XOR2_X1 U1096 ( .A(G286), .B(G171), .Z(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(n1013), .ZN(n1018) );
  XNOR2_X1 U1098 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(G37), .A2(n1019), .ZN(G397) );
  XOR2_X1 U1101 ( .A(G2446), .B(KEYINPUT106), .Z(n1021) );
  XNOR2_X1 U1102 ( .A(G2427), .B(G2443), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1021), .B(n1020), .ZN(n1022) );
  XOR2_X1 U1104 ( .A(n1022), .B(G2454), .Z(n1024) );
  XNOR2_X1 U1105 ( .A(G1348), .B(G2438), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(n1024), .B(n1023), .ZN(n1029) );
  XOR2_X1 U1107 ( .A(G2451), .B(KEYINPUT107), .Z(n1027) );
  XOR2_X1 U1108 ( .A(n1025), .B(G2435), .Z(n1026) );
  XNOR2_X1 U1109 ( .A(n1027), .B(n1026), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(n1029), .B(n1028), .Z(n1031) );
  XNOR2_X1 U1111 ( .A(KEYINPUT105), .B(G2430), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(n1031), .B(n1030), .ZN(n1032) );
  NAND2_X1 U1113 ( .A1(n1032), .A2(G14), .ZN(n1038) );
  NAND2_X1 U1114 ( .A1(G319), .A2(n1038), .ZN(n1035) );
  NOR2_X1 U1115 ( .A1(G227), .A2(G229), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(KEYINPUT49), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1037) );
  NOR2_X1 U1118 ( .A1(G395), .A2(G397), .ZN(n1036) );
  NAND2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(G225) );
  INV_X1 U1120 ( .A(G225), .ZN(G308) );
  INV_X1 U1121 ( .A(n1038), .ZN(G401) );
endmodule

