

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741;

  INV_X1 U371 ( .A(n649), .ZN(n645) );
  XOR2_X1 U372 ( .A(G122), .B(G107), .Z(n521) );
  XNOR2_X1 U373 ( .A(G143), .B(G113), .ZN(n507) );
  XNOR2_X1 U374 ( .A(G128), .B(G110), .ZN(n488) );
  XNOR2_X2 U375 ( .A(n572), .B(KEYINPUT1), .ZN(n663) );
  XNOR2_X2 U376 ( .A(n630), .B(n629), .ZN(n397) );
  XOR2_X2 U377 ( .A(n479), .B(KEYINPUT62), .Z(n409) );
  XOR2_X2 U378 ( .A(n694), .B(n693), .Z(n394) );
  NOR2_X2 U379 ( .A1(n561), .A2(n467), .ZN(n476) );
  XOR2_X2 U380 ( .A(n702), .B(KEYINPUT121), .Z(n704) );
  XNOR2_X2 U381 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X2 U382 ( .A(G902), .B(KEYINPUT15), .Z(n496) );
  XNOR2_X1 U383 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n361) );
  XNOR2_X1 U384 ( .A(G116), .B(G134), .ZN(n520) );
  INV_X1 U385 ( .A(G110), .ZN(n360) );
  INV_X2 U386 ( .A(KEYINPUT64), .ZN(n369) );
  INV_X1 U387 ( .A(n383), .ZN(n661) );
  AND2_X1 U388 ( .A1(n483), .A2(G224), .ZN(n348) );
  XNOR2_X1 U389 ( .A(KEYINPUT38), .B(n569), .ZN(n349) );
  NOR2_X2 U390 ( .A1(n740), .A2(n736), .ZN(n592) );
  NOR2_X1 U391 ( .A1(n641), .A2(n645), .ZN(n532) );
  NAND2_X1 U392 ( .A1(n387), .A2(n349), .ZN(n587) );
  NAND2_X2 U393 ( .A1(n657), .A2(n658), .ZN(n662) );
  XNOR2_X1 U394 ( .A(n360), .B(G107), .ZN(n707) );
  NAND2_X1 U395 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X2 U396 ( .A(G119), .B(KEYINPUT23), .ZN(n487) );
  INV_X2 U397 ( .A(G104), .ZN(n353) );
  INV_X1 U398 ( .A(KEYINPUT70), .ZN(n352) );
  INV_X1 U399 ( .A(G237), .ZN(n372) );
  INV_X1 U400 ( .A(G953), .ZN(n373) );
  NOR2_X1 U401 ( .A1(n739), .A2(KEYINPUT44), .ZN(n442) );
  XNOR2_X1 U402 ( .A(n589), .B(n588), .ZN(n736) );
  AND2_X1 U403 ( .A1(n645), .A2(n623), .ZN(n589) );
  BUF_X1 U404 ( .A(n556), .Z(n739) );
  XNOR2_X1 U405 ( .A(n587), .B(KEYINPUT39), .ZN(n623) );
  XNOR2_X1 U406 ( .A(n416), .B(n546), .ZN(n556) );
  XNOR2_X1 U407 ( .A(n581), .B(n580), .ZN(n740) );
  XNOR2_X1 U408 ( .A(n506), .B(n404), .ZN(n403) );
  OR2_X1 U409 ( .A1(n600), .A2(n685), .ZN(n581) );
  INV_X1 U410 ( .A(n594), .ZN(n387) );
  XNOR2_X1 U411 ( .A(n388), .B(KEYINPUT76), .ZN(n594) );
  AND2_X1 U412 ( .A1(n382), .A2(n661), .ZN(n381) );
  NOR2_X2 U413 ( .A1(n572), .A2(n662), .ZN(n584) );
  NOR2_X1 U414 ( .A1(n563), .A2(n586), .ZN(n573) );
  NAND2_X1 U415 ( .A1(n544), .A2(n542), .ZN(n649) );
  XNOR2_X1 U416 ( .A(n481), .B(n480), .ZN(n383) );
  XNOR2_X1 U417 ( .A(n518), .B(n519), .ZN(n544) );
  NOR2_X1 U418 ( .A1(G902), .A2(n479), .ZN(n481) );
  OR2_X1 U419 ( .A1(n697), .A2(G902), .ZN(n399) );
  XNOR2_X1 U420 ( .A(n462), .B(n384), .ZN(n479) );
  XNOR2_X1 U421 ( .A(n516), .B(n378), .ZN(n630) );
  XNOR2_X1 U422 ( .A(n380), .B(n379), .ZN(n378) );
  XNOR2_X1 U423 ( .A(n513), .B(n517), .ZN(n380) );
  XNOR2_X1 U424 ( .A(n355), .B(n469), .ZN(n708) );
  XNOR2_X1 U425 ( .A(n460), .B(n386), .ZN(n385) );
  XNOR2_X1 U426 ( .A(n370), .B(n348), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n470), .B(KEYINPUT16), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n515), .B(n352), .ZN(n470) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n489) );
  INV_X1 U430 ( .A(n707), .ZN(n359) );
  XNOR2_X1 U431 ( .A(n371), .B(KEYINPUT75), .ZN(n509) );
  XNOR2_X1 U432 ( .A(n512), .B(KEYINPUT101), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n354), .B(n358), .ZN(n469) );
  XNOR2_X1 U434 ( .A(n456), .B(KEYINPUT3), .ZN(n358) );
  XNOR2_X1 U435 ( .A(n487), .B(KEYINPUT93), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n461), .B(G137), .ZN(n386) );
  XNOR2_X1 U437 ( .A(n357), .B(n356), .ZN(n354) );
  XNOR2_X1 U438 ( .A(n353), .B(G122), .ZN(n515) );
  XNOR2_X2 U439 ( .A(G119), .B(KEYINPUT67), .ZN(n356) );
  INV_X2 U440 ( .A(KEYINPUT69), .ZN(n362) );
  XNOR2_X1 U441 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n510) );
  INV_X1 U442 ( .A(KEYINPUT90), .ZN(n456) );
  XNOR2_X1 U443 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n376) );
  XOR2_X2 U444 ( .A(G131), .B(G134), .Z(n723) );
  XNOR2_X2 U445 ( .A(G116), .B(G113), .ZN(n357) );
  XNOR2_X1 U446 ( .A(n350), .B(n359), .ZN(n364) );
  XNOR2_X1 U447 ( .A(n351), .B(n361), .ZN(n350) );
  XNOR2_X1 U448 ( .A(n351), .B(n707), .ZN(n468) );
  XNOR2_X2 U449 ( .A(n362), .B(KEYINPUT68), .ZN(n351) );
  XNOR2_X2 U450 ( .A(n459), .B(G143), .ZN(n523) );
  XNOR2_X1 U451 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U452 ( .A(n368), .B(n365), .ZN(n471) );
  XNOR2_X2 U453 ( .A(n725), .B(G101), .ZN(n368) );
  XNOR2_X2 U454 ( .A(n523), .B(KEYINPUT4), .ZN(n725) );
  XNOR2_X2 U455 ( .A(G125), .B(G146), .ZN(n367) );
  XNOR2_X1 U456 ( .A(n367), .B(n366), .ZN(n370) );
  INV_X1 U457 ( .A(KEYINPUT91), .ZN(n366) );
  XNOR2_X1 U458 ( .A(n367), .B(KEYINPUT10), .ZN(n514) );
  XNOR2_X2 U459 ( .A(n369), .B(G953), .ZN(n483) );
  XNOR2_X1 U460 ( .A(n368), .B(n385), .ZN(n384) );
  XNOR2_X1 U461 ( .A(n368), .B(n468), .ZN(n392) );
  NAND2_X1 U462 ( .A1(n374), .A2(n575), .ZN(n576) );
  XNOR2_X1 U463 ( .A(n375), .B(n574), .ZN(n374) );
  NAND2_X1 U464 ( .A1(n573), .A2(n383), .ZN(n375) );
  NAND2_X1 U465 ( .A1(n383), .A2(n671), .ZN(n583) );
  INV_X1 U466 ( .A(n657), .ZN(n382) );
  XNOR2_X1 U467 ( .A(n661), .B(KEYINPUT6), .ZN(n564) );
  AND2_X1 U468 ( .A1(n539), .A2(n383), .ZN(n668) );
  NAND2_X1 U469 ( .A1(n585), .A2(n389), .ZN(n388) );
  AND2_X1 U470 ( .A1(n584), .A2(n390), .ZN(n389) );
  INV_X1 U471 ( .A(n586), .ZN(n390) );
  BUF_X1 U472 ( .A(n688), .Z(n391) );
  XNOR2_X1 U473 ( .A(n549), .B(KEYINPUT85), .ZN(n443) );
  OR2_X2 U474 ( .A1(n429), .A2(n427), .ZN(n699) );
  XNOR2_X1 U475 ( .A(n393), .B(n394), .ZN(n695) );
  NOR2_X1 U476 ( .A1(n688), .A2(n424), .ZN(n393) );
  NOR2_X1 U477 ( .A1(n663), .A2(n662), .ZN(n539) );
  XOR2_X1 U478 ( .A(G137), .B(G140), .Z(n494) );
  XNOR2_X1 U479 ( .A(n540), .B(n396), .ZN(n414) );
  NAND2_X1 U480 ( .A1(n442), .A2(n441), .ZN(n440) );
  OR2_X1 U481 ( .A1(n625), .A2(n425), .ZN(n423) );
  INV_X1 U482 ( .A(G475), .ZN(n425) );
  NOR2_X1 U483 ( .A1(n490), .A2(G952), .ZN(n706) );
  XOR2_X1 U484 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n461) );
  XOR2_X1 U485 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n511) );
  NAND2_X1 U486 ( .A1(G234), .A2(G237), .ZN(n463) );
  OR2_X1 U487 ( .A1(G237), .A2(G902), .ZN(n474) );
  XNOR2_X1 U488 ( .A(n418), .B(KEYINPUT34), .ZN(n417) );
  XNOR2_X1 U489 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n491) );
  XOR2_X1 U490 ( .A(G140), .B(G131), .Z(n508) );
  NOR2_X1 U491 ( .A1(n679), .A2(n402), .ZN(n680) );
  INV_X1 U492 ( .A(n414), .ZN(n402) );
  NAND2_X1 U493 ( .A1(n624), .A2(n656), .ZN(n729) );
  NOR2_X1 U494 ( .A1(n735), .A2(n622), .ZN(n624) );
  INV_X1 U495 ( .A(KEYINPUT45), .ZN(n444) );
  INV_X1 U496 ( .A(KEYINPUT22), .ZN(n448) );
  INV_X1 U497 ( .A(KEYINPUT31), .ZN(n404) );
  INV_X1 U498 ( .A(KEYINPUT111), .ZN(n405) );
  OR2_X1 U499 ( .A1(n625), .A2(n480), .ZN(n422) );
  INV_X1 U500 ( .A(G217), .ZN(n426) );
  INV_X1 U501 ( .A(G478), .ZN(n428) );
  INV_X1 U502 ( .A(G469), .ZN(n427) );
  XNOR2_X1 U503 ( .A(n486), .B(n401), .ZN(n400) );
  INV_X1 U504 ( .A(n482), .ZN(n401) );
  NAND2_X1 U505 ( .A1(n496), .A2(G210), .ZN(n424) );
  XNOR2_X1 U506 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n552) );
  INV_X1 U507 ( .A(n403), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n412), .B(n397), .ZN(n631) );
  XOR2_X1 U509 ( .A(KEYINPUT66), .B(G469), .Z(n395) );
  XNOR2_X1 U510 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n396) );
  XNOR2_X2 U511 ( .A(n398), .B(n475), .ZN(n598) );
  NOR2_X1 U512 ( .A1(n614), .A2(n398), .ZN(n615) );
  XNOR2_X2 U513 ( .A(n431), .B(KEYINPUT87), .ZN(n398) );
  XNOR2_X2 U514 ( .A(n399), .B(n395), .ZN(n572) );
  XNOR2_X1 U515 ( .A(n392), .B(n400), .ZN(n697) );
  NOR2_X1 U516 ( .A1(n685), .A2(n402), .ZN(n686) );
  XNOR2_X1 U517 ( .A(n405), .B(n576), .ZN(n600) );
  BUF_X1 U518 ( .A(n692), .Z(n694) );
  BUF_X1 U519 ( .A(n554), .Z(n406) );
  XNOR2_X1 U520 ( .A(n553), .B(n552), .ZN(n407) );
  XNOR2_X1 U521 ( .A(n553), .B(n552), .ZN(n738) );
  XNOR2_X1 U522 ( .A(n408), .B(n409), .ZN(n626) );
  NOR2_X1 U523 ( .A1(n688), .A2(n422), .ZN(n408) );
  NOR2_X1 U524 ( .A1(n439), .A2(n437), .ZN(n436) );
  NOR2_X1 U525 ( .A1(n443), .A2(n446), .ZN(n439) );
  BUF_X1 U526 ( .A(n598), .Z(n599) );
  BUF_X1 U527 ( .A(n523), .Z(n410) );
  BUF_X1 U528 ( .A(n725), .Z(n411) );
  NAND2_X2 U529 ( .A1(n551), .A2(n550), .ZN(n553) );
  OR2_X2 U530 ( .A1(n429), .A2(n426), .ZN(n703) );
  NOR2_X1 U531 ( .A1(n688), .A2(n423), .ZN(n412) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n568) );
  XNOR2_X1 U533 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U534 ( .A1(n413), .A2(KEYINPUT84), .ZN(n438) );
  INV_X1 U535 ( .A(n555), .ZN(n413) );
  AND2_X1 U536 ( .A1(n541), .A2(n414), .ZN(n418) );
  XNOR2_X2 U537 ( .A(n478), .B(n477), .ZN(n541) );
  NOR2_X2 U538 ( .A1(n631), .A2(n706), .ZN(n632) );
  XNOR2_X1 U539 ( .A(n415), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U540 ( .A1(n695), .A2(n706), .ZN(n415) );
  NAND2_X1 U541 ( .A1(n417), .A2(n545), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n633), .A2(n419), .ZN(n538) );
  NAND2_X1 U543 ( .A1(n420), .A2(n604), .ZN(n419) );
  NAND2_X1 U544 ( .A1(n403), .A2(n636), .ZN(n420) );
  NAND2_X1 U545 ( .A1(n554), .A2(n537), .ZN(n633) );
  AND2_X2 U546 ( .A1(n433), .A2(n663), .ZN(n554) );
  XNOR2_X2 U547 ( .A(n536), .B(n448), .ZN(n433) );
  NAND2_X1 U548 ( .A1(n421), .A2(n496), .ZN(n429) );
  INV_X1 U549 ( .A(n688), .ZN(n421) );
  OR2_X1 U550 ( .A1(n429), .A2(n428), .ZN(n452) );
  NAND2_X1 U551 ( .A1(n436), .A2(n434), .ZN(n445) );
  NOR2_X2 U552 ( .A1(n626), .A2(n706), .ZN(n628) );
  XNOR2_X2 U553 ( .A(n430), .B(KEYINPUT2), .ZN(n688) );
  NOR2_X2 U554 ( .A1(n716), .A2(n729), .ZN(n430) );
  XNOR2_X2 U555 ( .A(n445), .B(n444), .ZN(n716) );
  NOR2_X2 U556 ( .A1(n568), .A2(n432), .ZN(n431) );
  INV_X1 U557 ( .A(n671), .ZN(n432) );
  AND2_X1 U558 ( .A1(n433), .A2(n447), .ZN(n551) );
  NAND2_X1 U559 ( .A1(n443), .A2(n435), .ZN(n434) );
  AND2_X1 U560 ( .A1(n555), .A2(n446), .ZN(n435) );
  NAND2_X1 U561 ( .A1(n438), .A2(n440), .ZN(n437) );
  INV_X1 U562 ( .A(n557), .ZN(n441) );
  INV_X1 U563 ( .A(KEYINPUT84), .ZN(n446) );
  INV_X1 U564 ( .A(n564), .ZN(n447) );
  AND2_X1 U565 ( .A1(n449), .A2(n641), .ZN(n653) );
  AND2_X1 U566 ( .A1(n449), .A2(n645), .ZN(n651) );
  NOR2_X1 U567 ( .A1(n450), .A2(n706), .ZN(G63) );
  XNOR2_X1 U568 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U569 ( .A(n701), .B(KEYINPUT120), .ZN(n451) );
  XOR2_X1 U570 ( .A(n499), .B(n498), .Z(n453) );
  AND2_X1 U571 ( .A1(G221), .A2(n524), .ZN(n454) );
  AND2_X1 U572 ( .A1(n619), .A2(n655), .ZN(n455) );
  INV_X1 U573 ( .A(KEYINPUT83), .ZN(n590) );
  XNOR2_X1 U574 ( .A(n590), .B(KEYINPUT46), .ZN(n591) );
  XNOR2_X1 U575 ( .A(n592), .B(n591), .ZN(n620) );
  INV_X1 U576 ( .A(KEYINPUT19), .ZN(n475) );
  XOR2_X1 U577 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n458) );
  XOR2_X1 U578 ( .A(G146), .B(n723), .Z(n482) );
  XNOR2_X1 U579 ( .A(n469), .B(n482), .ZN(n457) );
  XNOR2_X1 U580 ( .A(n458), .B(n457), .ZN(n462) );
  XNOR2_X2 U581 ( .A(G128), .B(KEYINPUT65), .ZN(n459) );
  NAND2_X1 U582 ( .A1(G210), .A2(n509), .ZN(n460) );
  XOR2_X1 U583 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n464) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U585 ( .A1(G952), .A2(n465), .ZN(n684) );
  NOR2_X1 U586 ( .A1(G953), .A2(n684), .ZN(n561) );
  NAND2_X1 U587 ( .A1(G902), .A2(n465), .ZN(n558) );
  INV_X1 U588 ( .A(G898), .ZN(n466) );
  NAND2_X1 U589 ( .A1(G953), .A2(n466), .ZN(n711) );
  NOR2_X1 U590 ( .A1(n558), .A2(n711), .ZN(n467) );
  XNOR2_X1 U591 ( .A(n471), .B(n708), .ZN(n692) );
  NOR2_X1 U592 ( .A1(n692), .A2(n496), .ZN(n473) );
  AND2_X1 U593 ( .A1(G210), .A2(n474), .ZN(n472) );
  NAND2_X1 U594 ( .A1(G214), .A2(n474), .ZN(n671) );
  NOR2_X2 U595 ( .A1(n598), .A2(n476), .ZN(n478) );
  XNOR2_X1 U596 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n477) );
  INV_X1 U597 ( .A(G472), .ZN(n480) );
  XOR2_X1 U598 ( .A(G104), .B(n494), .Z(n485) );
  BUF_X2 U599 ( .A(n483), .Z(n490) );
  NAND2_X1 U600 ( .A1(G227), .A2(n490), .ZN(n484) );
  XNOR2_X1 U601 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n489), .B(n488), .ZN(n493) );
  NAND2_X1 U603 ( .A1(n490), .A2(G234), .ZN(n492) );
  XNOR2_X1 U604 ( .A(n492), .B(n491), .ZN(n524) );
  XNOR2_X1 U605 ( .A(n493), .B(n454), .ZN(n495) );
  XOR2_X1 U606 ( .A(n494), .B(n514), .Z(n722) );
  XNOR2_X1 U607 ( .A(n495), .B(n722), .ZN(n702) );
  NOR2_X1 U608 ( .A1(G902), .A2(n702), .ZN(n502) );
  INV_X1 U609 ( .A(n496), .ZN(n625) );
  NAND2_X1 U610 ( .A1(G234), .A2(n625), .ZN(n497) );
  XNOR2_X1 U611 ( .A(KEYINPUT20), .B(n497), .ZN(n503) );
  NAND2_X1 U612 ( .A1(n503), .A2(G217), .ZN(n500) );
  XOR2_X1 U613 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n499) );
  XNOR2_X1 U614 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n498) );
  XNOR2_X1 U615 ( .A(n500), .B(n453), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n562) );
  INV_X2 U617 ( .A(n562), .ZN(n657) );
  NAND2_X1 U618 ( .A1(n503), .A2(G221), .ZN(n504) );
  XOR2_X1 U619 ( .A(KEYINPUT21), .B(n504), .Z(n658) );
  AND2_X1 U620 ( .A1(n661), .A2(n584), .ZN(n505) );
  NAND2_X1 U621 ( .A1(n541), .A2(n505), .ZN(n636) );
  NAND2_X1 U622 ( .A1(n668), .A2(n541), .ZN(n506) );
  XNOR2_X1 U623 ( .A(KEYINPUT13), .B(G475), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n508), .B(n507), .ZN(n517) );
  NAND2_X1 U625 ( .A1(G214), .A2(n509), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U627 ( .A(n515), .B(n514), .ZN(n516) );
  NOR2_X1 U628 ( .A1(G902), .A2(n630), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U630 ( .A(n410), .B(n522), .ZN(n530) );
  NAND2_X1 U631 ( .A1(n524), .A2(G217), .ZN(n528) );
  XOR2_X1 U632 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n526) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n525) );
  XNOR2_X1 U634 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U635 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U636 ( .A(n530), .B(n529), .ZN(n701) );
  NOR2_X1 U637 ( .A1(n701), .A2(G902), .ZN(n531) );
  XNOR2_X1 U638 ( .A(n531), .B(G478), .ZN(n542) );
  NOR2_X1 U639 ( .A1(n544), .A2(n542), .ZN(n641) );
  XNOR2_X1 U640 ( .A(n532), .B(KEYINPUT104), .ZN(n675) );
  INV_X1 U641 ( .A(n675), .ZN(n604) );
  INV_X1 U642 ( .A(n663), .ZN(n618) );
  INV_X1 U643 ( .A(n544), .ZN(n533) );
  NAND2_X1 U644 ( .A1(n533), .A2(n542), .ZN(n673) );
  INV_X1 U645 ( .A(n658), .ZN(n534) );
  NOR2_X1 U646 ( .A1(n673), .A2(n534), .ZN(n535) );
  NAND2_X1 U647 ( .A1(n541), .A2(n535), .ZN(n536) );
  NOR2_X1 U648 ( .A1(n562), .A2(n564), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n538), .B(KEYINPUT105), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n539), .A2(n564), .ZN(n540) );
  INV_X1 U651 ( .A(n542), .ZN(n543) );
  NAND2_X1 U652 ( .A1(n544), .A2(n543), .ZN(n593) );
  XNOR2_X1 U653 ( .A(n593), .B(KEYINPUT77), .ZN(n545) );
  XNOR2_X1 U654 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n546) );
  NAND2_X1 U655 ( .A1(n556), .A2(KEYINPUT44), .ZN(n547) );
  NAND2_X1 U656 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U657 ( .A1(n663), .A2(n657), .ZN(n550) );
  NAND2_X1 U658 ( .A1(n406), .A2(n381), .ZN(n640) );
  NAND2_X1 U659 ( .A1(n738), .A2(n640), .ZN(n557) );
  NAND2_X1 U660 ( .A1(n557), .A2(KEYINPUT44), .ZN(n555) );
  OR2_X1 U661 ( .A1(n490), .A2(n558), .ZN(n559) );
  NOR2_X1 U662 ( .A1(G900), .A2(n559), .ZN(n560) );
  NOR2_X1 U663 ( .A1(n561), .A2(n560), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n562), .A2(n658), .ZN(n563) );
  AND2_X1 U665 ( .A1(n564), .A2(n645), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n573), .A2(n565), .ZN(n614) );
  NOR2_X1 U667 ( .A1(n618), .A2(n614), .ZN(n566) );
  NAND2_X1 U668 ( .A1(n566), .A2(n671), .ZN(n567) );
  XNOR2_X1 U669 ( .A(n567), .B(KEYINPUT43), .ZN(n570) );
  BUF_X1 U670 ( .A(n568), .Z(n569) );
  NAND2_X1 U671 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U672 ( .A(KEYINPUT107), .B(n571), .ZN(n735) );
  XNOR2_X1 U673 ( .A(n572), .B(KEYINPUT109), .ZN(n575) );
  XOR2_X1 U674 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n574) );
  NAND2_X1 U675 ( .A1(n349), .A2(n671), .ZN(n676) );
  NOR2_X1 U676 ( .A1(n676), .A2(n673), .ZN(n578) );
  XNOR2_X1 U677 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n577) );
  XOR2_X1 U678 ( .A(n578), .B(n577), .Z(n685) );
  XNOR2_X1 U679 ( .A(KEYINPUT42), .B(KEYINPUT114), .ZN(n579) );
  XNOR2_X1 U680 ( .A(n579), .B(KEYINPUT115), .ZN(n580) );
  XOR2_X1 U681 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n582) );
  XNOR2_X1 U682 ( .A(n583), .B(n582), .ZN(n585) );
  XNOR2_X1 U683 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n588) );
  INV_X1 U684 ( .A(n569), .ZN(n596) );
  NOR2_X1 U685 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n596), .A2(n595), .ZN(n644) );
  XNOR2_X1 U687 ( .A(KEYINPUT80), .B(n644), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n675), .A2(KEYINPUT47), .ZN(n597) );
  XOR2_X1 U689 ( .A(n597), .B(KEYINPUT79), .Z(n603) );
  NOR2_X2 U690 ( .A1(n600), .A2(n599), .ZN(n646) );
  NAND2_X1 U691 ( .A1(KEYINPUT72), .A2(n646), .ZN(n601) );
  NAND2_X1 U692 ( .A1(n601), .A2(KEYINPUT47), .ZN(n602) );
  NAND2_X1 U693 ( .A1(n603), .A2(n602), .ZN(n610) );
  INV_X1 U694 ( .A(n646), .ZN(n608) );
  XNOR2_X1 U695 ( .A(n604), .B(KEYINPUT72), .ZN(n606) );
  INV_X1 U696 ( .A(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U697 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U698 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U699 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U701 ( .A(n613), .B(KEYINPUT71), .ZN(n619) );
  XOR2_X1 U702 ( .A(KEYINPUT36), .B(KEYINPUT86), .Z(n616) );
  XOR2_X1 U703 ( .A(n616), .B(n615), .Z(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n655) );
  NAND2_X1 U705 ( .A1(n620), .A2(n455), .ZN(n621) );
  XNOR2_X1 U706 ( .A(n621), .B(KEYINPUT48), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n641), .ZN(n656) );
  XNOR2_X1 U708 ( .A(KEYINPUT63), .B(KEYINPUT89), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n628), .B(n627), .ZN(G57) );
  XOR2_X1 U710 ( .A(KEYINPUT119), .B(KEYINPUT59), .Z(n629) );
  XNOR2_X1 U711 ( .A(n632), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U712 ( .A(n633), .Z(n634) );
  XNOR2_X1 U713 ( .A(G101), .B(n634), .ZN(G3) );
  NOR2_X1 U714 ( .A1(n649), .A2(n636), .ZN(n635) );
  XOR2_X1 U715 ( .A(G104), .B(n635), .Z(G6) );
  INV_X1 U716 ( .A(n641), .ZN(n652) );
  NOR2_X1 U717 ( .A1(n652), .A2(n636), .ZN(n638) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U720 ( .A(G107), .B(n639), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(n640), .ZN(G12) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n643) );
  NAND2_X1 U723 ( .A1(n646), .A2(n641), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n643), .B(n642), .ZN(G30) );
  XNOR2_X1 U725 ( .A(G143), .B(n644), .ZN(G45) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n647), .B(KEYINPUT116), .ZN(n648) );
  XNOR2_X1 U728 ( .A(G146), .B(n648), .ZN(G48) );
  XNOR2_X1 U729 ( .A(G113), .B(KEYINPUT117), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n651), .B(n650), .ZN(G15) );
  XOR2_X1 U731 ( .A(G116), .B(n653), .Z(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n656), .ZN(G36) );
  NOR2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(KEYINPUT49), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n666) );
  AND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(KEYINPUT50), .ZN(n665) );
  NOR2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT51), .B(n669), .Z(n670) );
  NOR2_X1 U743 ( .A1(n685), .A2(n670), .ZN(n681) );
  NOR2_X1 U744 ( .A1(n349), .A2(n671), .ZN(n672) );
  NOR2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U746 ( .A(n674), .B(KEYINPUT118), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n689), .A2(n391), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n690), .A2(G953), .ZN(n691) );
  XNOR2_X1 U755 ( .A(n691), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U756 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n693) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  NOR2_X1 U758 ( .A1(n706), .A2(n700), .ZN(G54) );
  XNOR2_X1 U759 ( .A(n703), .B(n704), .ZN(n705) );
  NOR2_X1 U760 ( .A1(n706), .A2(n705), .ZN(G66) );
  XNOR2_X1 U761 ( .A(G101), .B(n707), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n721) );
  NAND2_X1 U764 ( .A1(G224), .A2(G953), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(KEYINPUT61), .ZN(n713) );
  XNOR2_X1 U766 ( .A(KEYINPUT122), .B(n713), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n714), .A2(G898), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT123), .ZN(n719) );
  BUF_X1 U769 ( .A(n716), .Z(n717) );
  NOR2_X1 U770 ( .A1(n717), .A2(G953), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(G69) );
  XOR2_X1 U773 ( .A(n723), .B(n722), .Z(n724) );
  XNOR2_X1 U774 ( .A(n411), .B(n724), .ZN(n730) );
  XNOR2_X1 U775 ( .A(G227), .B(n730), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G900), .ZN(n727) );
  XNOR2_X1 U777 ( .A(KEYINPUT124), .B(n727), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n728), .A2(G953), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(n490), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(n734), .Z(G72) );
  XOR2_X1 U783 ( .A(G140), .B(n735), .Z(G42) );
  XNOR2_X1 U784 ( .A(G131), .B(n736), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n737), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U786 ( .A(n407), .B(G119), .ZN(G21) );
  XOR2_X1 U787 ( .A(n739), .B(G122), .Z(G24) );
  XOR2_X1 U788 ( .A(G137), .B(n740), .Z(n741) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n741), .ZN(G39) );
endmodule

