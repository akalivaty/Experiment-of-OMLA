

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600;

  XNOR2_X1 U324 ( .A(n375), .B(n374), .ZN(n376) );
  NAND2_X1 U325 ( .A1(n454), .A2(n594), .ZN(n455) );
  NOR2_X1 U326 ( .A1(n481), .A2(n534), .ZN(n483) );
  XNOR2_X1 U327 ( .A(n490), .B(KEYINPUT37), .ZN(n513) );
  NAND2_X1 U328 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U329 ( .A(n385), .B(n384), .Z(n526) );
  XNOR2_X1 U330 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U331 ( .A(G43GAT), .B(KEYINPUT7), .Z(n292) );
  AND2_X1 U332 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U333 ( .A(KEYINPUT40), .B(n519), .Z(n294) );
  INV_X1 U334 ( .A(KEYINPUT45), .ZN(n451) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U336 ( .A(n461), .B(KEYINPUT119), .ZN(n462) );
  INV_X1 U337 ( .A(KEYINPUT103), .ZN(n482) );
  XNOR2_X1 U338 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U339 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U340 ( .A(G8GAT), .B(G169GAT), .Z(n409) );
  NOR2_X1 U341 ( .A1(n534), .A2(n464), .ZN(n465) );
  NOR2_X1 U342 ( .A1(n457), .A2(n456), .ZN(n459) );
  INV_X1 U343 ( .A(KEYINPUT100), .ZN(n374) );
  OR2_X1 U344 ( .A1(n543), .A2(n567), .ZN(n349) );
  XNOR2_X1 U345 ( .A(n389), .B(n293), .ZN(n340) );
  XNOR2_X1 U346 ( .A(n349), .B(KEYINPUT26), .ZN(n475) );
  XNOR2_X1 U347 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U348 ( .A(n341), .B(n340), .ZN(n348) );
  NOR2_X1 U349 ( .A1(n475), .A2(n466), .ZN(n587) );
  XNOR2_X1 U350 ( .A(n406), .B(n405), .ZN(n453) );
  INV_X1 U351 ( .A(KEYINPUT126), .ZN(n468) );
  XNOR2_X1 U352 ( .A(n491), .B(KEYINPUT111), .ZN(n539) );
  XNOR2_X1 U353 ( .A(n515), .B(KEYINPUT38), .ZN(n520) );
  XNOR2_X1 U354 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U355 ( .A(n493), .B(n295), .ZN(n494) );
  XNOR2_X1 U356 ( .A(n471), .B(n470), .ZN(G1355GAT) );
  XNOR2_X1 U357 ( .A(n495), .B(n494), .ZN(G1339GAT) );
  INV_X1 U358 ( .A(G106GAT), .ZN(n295) );
  XOR2_X1 U359 ( .A(G92GAT), .B(G106GAT), .Z(n297) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n296) );
  XNOR2_X1 U361 ( .A(n297), .B(n296), .ZN(n312) );
  XOR2_X1 U362 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n299) );
  NAND2_X1 U363 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U364 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U365 ( .A(n300), .B(KEYINPUT66), .Z(n304) );
  XNOR2_X1 U366 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n301) );
  XNOR2_X1 U367 ( .A(n301), .B(G99GAT), .ZN(n399) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U369 ( .A(n292), .B(n302), .ZN(n418) );
  XNOR2_X1 U370 ( .A(n399), .B(n418), .ZN(n303) );
  XNOR2_X1 U371 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U372 ( .A(KEYINPUT11), .B(KEYINPUT79), .Z(n306) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n305) );
  XNOR2_X1 U374 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U375 ( .A(n308), .B(n307), .Z(n310) );
  XOR2_X1 U376 ( .A(G190GAT), .B(G36GAT), .Z(n373) );
  XOR2_X1 U377 ( .A(G162GAT), .B(G50GAT), .Z(n334) );
  XNOR2_X1 U378 ( .A(n373), .B(n334), .ZN(n309) );
  XNOR2_X1 U379 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X2 U380 ( .A(n312), .B(n311), .Z(n583) );
  XNOR2_X1 U381 ( .A(KEYINPUT36), .B(n583), .ZN(n488) );
  XOR2_X1 U382 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n314) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(KEYINPUT89), .ZN(n313) );
  XNOR2_X1 U384 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U385 ( .A(G127GAT), .B(G15GAT), .Z(n436) );
  XOR2_X1 U386 ( .A(n315), .B(n436), .Z(n317) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U388 ( .A(n317), .B(n316), .ZN(n323) );
  XOR2_X1 U389 ( .A(G113GAT), .B(KEYINPUT0), .Z(n319) );
  XNOR2_X1 U390 ( .A(G134GAT), .B(KEYINPUT85), .ZN(n318) );
  XNOR2_X1 U391 ( .A(n319), .B(n318), .ZN(n363) );
  XOR2_X1 U392 ( .A(G120GAT), .B(G71GAT), .Z(n387) );
  XOR2_X1 U393 ( .A(n363), .B(n387), .Z(n321) );
  NAND2_X1 U394 ( .A1(G227GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U395 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U396 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U397 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n325) );
  XNOR2_X1 U398 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n324) );
  XNOR2_X1 U399 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U400 ( .A(G183GAT), .B(n326), .Z(n383) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G176GAT), .Z(n328) );
  XNOR2_X1 U402 ( .A(KEYINPUT87), .B(KEYINPUT90), .ZN(n327) );
  XNOR2_X1 U403 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U404 ( .A(n383), .B(n329), .ZN(n330) );
  XOR2_X1 U405 ( .A(n331), .B(n330), .Z(n507) );
  INV_X1 U406 ( .A(n507), .ZN(n543) );
  XOR2_X1 U407 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n333) );
  XNOR2_X1 U408 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n332) );
  XNOR2_X1 U409 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U410 ( .A(G155GAT), .B(G22GAT), .Z(n437) );
  XNOR2_X1 U411 ( .A(n334), .B(n437), .ZN(n336) );
  XOR2_X1 U412 ( .A(KEYINPUT22), .B(G204GAT), .Z(n335) );
  XNOR2_X1 U413 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U414 ( .A(n338), .B(n337), .Z(n341) );
  XNOR2_X1 U415 ( .A(G148GAT), .B(G106GAT), .ZN(n339) );
  XNOR2_X1 U416 ( .A(n339), .B(G78GAT), .ZN(n389) );
  INV_X1 U417 ( .A(n389), .ZN(n386) );
  XOR2_X1 U418 ( .A(G141GAT), .B(KEYINPUT3), .Z(n343) );
  XNOR2_X1 U419 ( .A(KEYINPUT94), .B(KEYINPUT2), .ZN(n342) );
  XNOR2_X1 U420 ( .A(n343), .B(n342), .ZN(n352) );
  XOR2_X1 U421 ( .A(KEYINPUT93), .B(G197GAT), .Z(n345) );
  XNOR2_X1 U422 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n344) );
  XNOR2_X1 U423 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U424 ( .A(G211GAT), .B(n346), .Z(n382) );
  XNOR2_X1 U425 ( .A(n352), .B(n382), .ZN(n347) );
  XNOR2_X1 U426 ( .A(n348), .B(n347), .ZN(n567) );
  XOR2_X1 U427 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n351) );
  XNOR2_X1 U428 ( .A(KEYINPUT4), .B(KEYINPUT95), .ZN(n350) );
  XNOR2_X1 U429 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U430 ( .A(n352), .B(KEYINPUT96), .Z(n354) );
  NAND2_X1 U431 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U432 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U433 ( .A(n356), .B(n355), .ZN(n370) );
  XOR2_X1 U434 ( .A(G57GAT), .B(G127GAT), .Z(n358) );
  XNOR2_X1 U435 ( .A(G155GAT), .B(G120GAT), .ZN(n357) );
  XNOR2_X1 U436 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U437 ( .A(KEYINPUT98), .B(KEYINPUT6), .Z(n360) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n359) );
  XNOR2_X1 U439 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U440 ( .A(n362), .B(n361), .Z(n368) );
  XOR2_X1 U441 ( .A(G85GAT), .B(G162GAT), .Z(n365) );
  XNOR2_X1 U442 ( .A(G148GAT), .B(n363), .ZN(n364) );
  XNOR2_X1 U443 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U444 ( .A(G29GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U445 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U446 ( .A(n370), .B(n369), .Z(n534) );
  XOR2_X1 U447 ( .A(n409), .B(KEYINPUT101), .Z(n372) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U449 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n373), .B(KEYINPUT99), .ZN(n375) );
  XOR2_X1 U451 ( .A(G204GAT), .B(KEYINPUT76), .Z(n379) );
  XNOR2_X1 U452 ( .A(G92GAT), .B(G176GAT), .ZN(n378) );
  XNOR2_X1 U453 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U454 ( .A(G64GAT), .B(n380), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n381), .B(n404), .ZN(n385) );
  XNOR2_X1 U456 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U457 ( .A(n526), .B(KEYINPUT118), .Z(n460) );
  NAND2_X1 U458 ( .A1(n386), .A2(n387), .ZN(n391) );
  INV_X1 U459 ( .A(n387), .ZN(n388) );
  NAND2_X1 U460 ( .A1(n389), .A2(n388), .ZN(n390) );
  NAND2_X1 U461 ( .A1(n391), .A2(n390), .ZN(n393) );
  NAND2_X1 U462 ( .A1(G230GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n396) );
  INV_X1 U464 ( .A(n396), .ZN(n394) );
  NAND2_X1 U465 ( .A1(n394), .A2(KEYINPUT32), .ZN(n398) );
  INV_X1 U466 ( .A(KEYINPUT32), .ZN(n395) );
  NAND2_X1 U467 ( .A1(n396), .A2(n395), .ZN(n397) );
  NAND2_X1 U468 ( .A1(n398), .A2(n397), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n399), .B(KEYINPUT33), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n402), .B(KEYINPUT74), .ZN(n406) );
  XOR2_X1 U472 ( .A(G57GAT), .B(KEYINPUT13), .Z(n431) );
  XOR2_X1 U473 ( .A(n431), .B(KEYINPUT31), .Z(n403) );
  XNOR2_X1 U474 ( .A(n453), .B(KEYINPUT41), .ZN(n575) );
  INV_X1 U475 ( .A(n575), .ZN(n472) );
  XOR2_X1 U476 ( .A(G197GAT), .B(G50GAT), .Z(n408) );
  XNOR2_X1 U477 ( .A(G113GAT), .B(G36GAT), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U479 ( .A(n410), .B(n409), .Z(n412) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(G22GAT), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U482 ( .A(KEYINPUT70), .B(KEYINPUT73), .Z(n414) );
  XNOR2_X1 U483 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U485 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n417), .B(KEYINPUT72), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n418), .B(n434), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n422) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U492 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U493 ( .A(KEYINPUT69), .B(n423), .Z(n424) );
  XOR2_X1 U494 ( .A(n425), .B(n424), .Z(n588) );
  NOR2_X1 U495 ( .A1(n472), .A2(n588), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n426), .B(KEYINPUT46), .ZN(n427) );
  NOR2_X1 U497 ( .A1(n427), .A2(n583), .ZN(n449) );
  XOR2_X1 U498 ( .A(G64GAT), .B(G8GAT), .Z(n429) );
  XNOR2_X1 U499 ( .A(G71GAT), .B(G183GAT), .ZN(n428) );
  XNOR2_X1 U500 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U501 ( .A(n430), .B(G211GAT), .Z(n433) );
  XNOR2_X1 U502 ( .A(n431), .B(G78GAT), .ZN(n432) );
  XNOR2_X1 U503 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U504 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U505 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U507 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n441) );
  NAND2_X1 U508 ( .A1(G231GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U509 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U510 ( .A(n443), .B(n442), .Z(n448) );
  XOR2_X1 U511 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n445) );
  XNOR2_X1 U512 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n444) );
  XNOR2_X1 U513 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U514 ( .A(n446), .B(KEYINPUT81), .ZN(n447) );
  XOR2_X1 U515 ( .A(n448), .B(n447), .Z(n580) );
  INV_X1 U516 ( .A(n580), .ZN(n598) );
  NAND2_X1 U517 ( .A1(n449), .A2(n598), .ZN(n450) );
  XNOR2_X1 U518 ( .A(n450), .B(KEYINPUT47), .ZN(n457) );
  INV_X1 U519 ( .A(n588), .ZN(n573) );
  NAND2_X1 U520 ( .A1(n488), .A2(n580), .ZN(n452) );
  BUF_X1 U521 ( .A(n453), .Z(n594) );
  NOR2_X1 U522 ( .A1(n573), .A2(n455), .ZN(n456) );
  INV_X1 U523 ( .A(KEYINPUT48), .ZN(n458) );
  XNOR2_X1 U524 ( .A(n459), .B(n458), .ZN(n542) );
  NAND2_X1 U525 ( .A1(n460), .A2(n542), .ZN(n463) );
  INV_X1 U526 ( .A(KEYINPUT54), .ZN(n461) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT64), .ZN(n568) );
  INV_X1 U528 ( .A(n568), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n488), .A2(n587), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(KEYINPUT62), .ZN(n471) );
  XNOR2_X1 U531 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n469) );
  NOR2_X1 U532 ( .A1(n472), .A2(n573), .ZN(n523) );
  XNOR2_X1 U533 ( .A(n526), .B(KEYINPUT27), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n473) );
  XOR2_X1 U535 ( .A(n567), .B(n473), .Z(n530) );
  INV_X1 U536 ( .A(n530), .ZN(n492) );
  NOR2_X1 U537 ( .A1(n476), .A2(n492), .ZN(n474) );
  NAND2_X1 U538 ( .A1(n474), .A2(n534), .ZN(n545) );
  NOR2_X1 U539 ( .A1(n543), .A2(n545), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n476), .A2(n475), .ZN(n555) );
  INV_X1 U541 ( .A(n526), .ZN(n536) );
  NAND2_X1 U542 ( .A1(n536), .A2(n543), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n477), .A2(n567), .ZN(n479) );
  XNOR2_X1 U544 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n478) );
  XNOR2_X1 U545 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U546 ( .A1(n555), .A2(n480), .ZN(n481) );
  NOR2_X1 U547 ( .A1(n485), .A2(n484), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(n486), .Z(n499) );
  NAND2_X1 U549 ( .A1(n598), .A2(n499), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(KEYINPUT109), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n523), .A2(n513), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n539), .A2(n492), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n493) );
  INV_X1 U554 ( .A(n534), .ZN(n557) );
  NAND2_X1 U555 ( .A1(n594), .A2(n573), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT77), .ZN(n514) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n498) );
  NOR2_X1 U558 ( .A1(n583), .A2(n598), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT105), .ZN(n522) );
  NAND2_X1 U562 ( .A1(n514), .A2(n522), .ZN(n510) );
  NOR2_X1 U563 ( .A1(n557), .A2(n510), .ZN(n503) );
  XNOR2_X1 U564 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U566 ( .A(G1GAT), .B(n504), .Z(G1324GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n510), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1325GAT) );
  BUF_X1 U570 ( .A(n507), .Z(n572) );
  NOR2_X1 U571 ( .A1(n572), .A2(n510), .ZN(n509) );
  XNOR2_X1 U572 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NOR2_X1 U574 ( .A1(n530), .A2(n510), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n515) );
  NOR2_X1 U578 ( .A1(n520), .A2(n557), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(KEYINPUT39), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G29GAT), .B(n517), .ZN(G1328GAT) );
  NOR2_X1 U581 ( .A1(n520), .A2(n526), .ZN(n518) );
  XOR2_X1 U582 ( .A(G36GAT), .B(n518), .Z(G1329GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n572), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G43GAT), .B(n294), .ZN(G1330GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n530), .ZN(n521) );
  XOR2_X1 U586 ( .A(G50GAT), .B(n521), .Z(G1331GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n557), .A2(n529), .ZN(n524) );
  XOR2_X1 U589 ( .A(G57GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT42), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n529), .ZN(n527) );
  XOR2_X1 U592 ( .A(G64GAT), .B(n527), .Z(G1333GAT) );
  NOR2_X1 U593 ( .A1(n572), .A2(n529), .ZN(n528) );
  XOR2_X1 U594 ( .A(G71GAT), .B(n528), .Z(G1334GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G78GAT), .B(n533), .ZN(G1335GAT) );
  NAND2_X1 U599 ( .A1(n539), .A2(n534), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U601 ( .A1(n539), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT112), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G92GAT), .B(n538), .ZN(G1337GAT) );
  XOR2_X1 U604 ( .A(G99GAT), .B(KEYINPUT113), .Z(n541) );
  NAND2_X1 U605 ( .A1(n539), .A2(n543), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1338GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n573), .A2(n551), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U612 ( .A1(n551), .A2(n575), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  NAND2_X1 U614 ( .A1(n580), .A2(n551), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(KEYINPUT50), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n583), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(G134GAT), .B(n554), .Z(G1343GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n542), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n573), .A2(n564), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n560) );
  NAND2_X1 U626 ( .A1(n564), .A2(n575), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n561), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n580), .A2(n564), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT116), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G155GAT), .B(n563), .ZN(G1346GAT) );
  XOR2_X1 U632 ( .A(G162GAT), .B(KEYINPUT117), .Z(n566) );
  NAND2_X1 U633 ( .A1(n564), .A2(n583), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n570) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  NOR2_X2 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G169GAT), .B(n574), .ZN(G1348GAT) );
  NAND2_X1 U641 ( .A1(n584), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G176GAT), .B(KEYINPUT57), .Z(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1349GAT) );
  NAND2_X1 U646 ( .A1(n580), .A2(n584), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT122), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(KEYINPUT58), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G190GAT), .B(n586), .ZN(G1351GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n597) );
  NOR2_X1 U653 ( .A1(n588), .A2(n597), .ZN(n593) );
  XOR2_X1 U654 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n590) );
  XNOR2_X1 U655 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(KEYINPUT60), .B(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1352GAT) );
  NOR2_X1 U659 ( .A1(n594), .A2(n597), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n596), .B(n595), .ZN(G1353GAT) );
  NOR2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U663 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n600), .B(n599), .ZN(G1354GAT) );
endmodule

