//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965;
  AND2_X1   g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G155gat), .B(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n210), .B2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n213), .B(new_n204), .C1(new_n212), .C2(new_n207), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT81), .B(G162gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G155gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n203), .B1(new_n218), .B2(KEYINPUT3), .ZN(new_n219));
  XNOR2_X1  g018(.A(G211gat), .B(G218gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G211gat), .A2(G218gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n220), .A2(new_n224), .A3(new_n223), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT29), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n218), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n227), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(new_n225), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n234));
  OAI211_X1 g033(.A(new_n211), .B(new_n234), .C1(new_n214), .C2(new_n217), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT85), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n232), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT85), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n229), .A4(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n218), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n236), .B1(new_n231), .B2(new_n225), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(KEYINPUT84), .ZN(new_n246));
  INV_X1    g045(.A(new_n234), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n245), .B2(KEYINPUT84), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n203), .B1(new_n249), .B2(new_n237), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n243), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g053(.A(G78gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n243), .A2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(G78gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n252), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT31), .B(G50gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G106gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n255), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n255), .B2(new_n259), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n267), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT70), .B1(new_n268), .B2(new_n267), .ZN(new_n270));
  OAI221_X1 g069(.A(new_n266), .B1(new_n267), .B2(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT27), .B(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n273), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n280));
  OAI211_X1 g079(.A(new_n271), .B(new_n279), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n266), .A2(KEYINPUT23), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n275), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n290), .B(new_n291), .C1(new_n273), .C2(KEYINPUT24), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n285), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n288), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n272), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n272), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n307), .A2(new_n308), .B1(new_n289), .B2(new_n275), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n298), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n295), .B1(new_n310), .B2(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n290), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n302), .B2(new_n304), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n314), .A2(new_n315), .A3(new_n298), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n281), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G127gat), .B(G134gat), .Z(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT1), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT72), .B(G120gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n323), .ZN(new_n327));
  XNOR2_X1  g126(.A(G113gat), .B(G120gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT1), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n329), .B2(new_n328), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n326), .A2(new_n327), .B1(new_n318), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G227gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n318), .ZN(new_n337));
  INV_X1    g136(.A(new_n327), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT73), .B1(new_n319), .B2(new_n323), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n281), .C1(new_n311), .C2(new_n316), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n342), .A2(KEYINPUT32), .ZN(new_n343));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT33), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n342), .B2(KEYINPUT32), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n343), .A2(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT34), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n341), .ZN(new_n356));
  INV_X1    g155(.A(new_n336), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT34), .B(new_n336), .C1(new_n333), .C2(new_n341), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n265), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n353), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n342), .A2(KEYINPUT32), .A3(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n360), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n360), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n264), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n340), .B2(new_n218), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n332), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n340), .A2(new_n235), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT83), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n332), .A2(new_n244), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n340), .A2(new_n218), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n378), .A2(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n374), .A2(new_n377), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(KEYINPUT5), .A3(new_n381), .A4(new_n375), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G1gat), .B(G29gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(G57gat), .B(G85gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395));
  INV_X1    g194(.A(new_n393), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n386), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n388), .A4(new_n396), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n315), .B1(new_n314), .B2(new_n298), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n295), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n281), .ZN(new_n406));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n401), .A2(KEYINPUT79), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n408), .A3(new_n406), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n404), .B2(new_n281), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n233), .B(new_n409), .C1(new_n410), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n406), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n408), .A3(new_n281), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n232), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n414), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT30), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n418), .B1(new_n414), .B2(new_n423), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n417), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n400), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT35), .B1(new_n372), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n398), .A2(new_n399), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n417), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n424), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n369), .A2(new_n370), .B1(new_n365), .B2(new_n364), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n264), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT40), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n382), .A2(new_n383), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n443), .B2(new_n380), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n380), .B2(new_n378), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n378), .A2(new_n446), .A3(new_n380), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n393), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n442), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n397), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n445), .A2(new_n448), .A3(new_n442), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n430), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n264), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n435), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n428), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n417), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n232), .B(new_n409), .C1(new_n410), .C2(new_n413), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n232), .B1(new_n420), .B2(new_n421), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n464), .A2(new_n463), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n455), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n414), .A2(KEYINPUT37), .A3(new_n423), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n459), .B1(new_n428), .B2(new_n456), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT87), .B(KEYINPUT37), .C1(new_n414), .C2(new_n423), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n418), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT38), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n454), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT76), .B1(new_n354), .B2(new_n360), .ZN(new_n477));
  AND4_X1   g276(.A1(KEYINPUT76), .A2(new_n360), .A3(new_n362), .A4(new_n363), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n477), .A2(new_n478), .B1(new_n360), .B2(new_n354), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n264), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n432), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n441), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488));
  INV_X1    g287(.A(G57gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n488), .B(G64gat), .C1(new_n489), .C2(KEYINPUT94), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n491));
  INV_X1    g290(.A(G64gat), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n491), .B(G57gat), .C1(new_n492), .C2(KEYINPUT93), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT93), .B1(new_n492), .B2(G57gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G71gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n258), .ZN(new_n497));
  NAND2_X1  g296(.A1(G71gat), .A2(G78gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n497), .A2(KEYINPUT95), .A3(new_n498), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n495), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n498), .B(new_n497), .C1(new_n506), .C2(new_n503), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT21), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT96), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT91), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AND4_X1   g321(.A1(new_n515), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n517), .A2(new_n518), .B1(new_n521), .B2(new_n516), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n515), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n507), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT97), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(KEYINPUT97), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n529), .B(KEYINPUT97), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n512), .A3(new_n513), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G183gat), .B(G211gat), .Z(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n532), .A2(new_n534), .A3(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  AND2_X1   g344(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT89), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G43gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G50gat), .ZN(new_n553));
  INV_X1    g352(.A(G50gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G43gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT15), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n551), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n550), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n553), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n555), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n559), .B(new_n560), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n558), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT14), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n549), .ZN(new_n569));
  NAND2_X1  g368(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n570));
  AOI21_X1  g369(.A(G36gat), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n550), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n567), .B(new_n556), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n556), .B1(new_n559), .B2(new_n567), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n565), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT17), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT98), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(G99gat), .A3(G106gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n581), .A3(KEYINPUT8), .ZN(new_n582));
  OR2_X1    g381(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(G85gat), .A3(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n582), .A2(new_n586), .A3(new_n591), .A4(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n566), .A2(new_n577), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n566), .A2(new_n577), .A3(new_n600), .A4(new_n597), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(new_n576), .B2(new_n597), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n599), .B(new_n601), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI22_X1  g413(.A1(new_n609), .A2(new_n610), .B1(KEYINPUT102), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n607), .A2(new_n608), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n608), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n613), .B(KEYINPUT102), .Z(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n566), .A2(new_n577), .A3(new_n526), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n557), .B(new_n565), .C1(new_n523), .C2(new_n525), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n621), .A2(KEYINPUT18), .A3(new_n622), .A4(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n526), .A2(new_n576), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(KEYINPUT92), .A3(new_n623), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n622), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n526), .A2(new_n631), .A3(new_n576), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G197gat), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT11), .B(G169gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n633), .A3(new_n640), .A4(new_n627), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT104), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n595), .A2(new_n505), .A3(new_n596), .A4(new_n507), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT103), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n597), .A2(new_n528), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(KEYINPUT103), .A3(KEYINPUT10), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n650), .ZN(new_n658));
  INV_X1    g457(.A(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n649), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n660), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n664), .B2(new_n648), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n657), .A2(new_n660), .A3(new_n666), .A4(new_n649), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n662), .A2(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR4_X1   g468(.A1(new_n544), .A2(new_n620), .A3(new_n644), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n487), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n400), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(new_n518), .ZN(G1324gat));
  INV_X1    g472(.A(new_n671), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n427), .A2(new_n431), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT107), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(G8gat), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(G1325gat));
  OR3_X1    g481(.A1(new_n671), .A2(G15gat), .A3(new_n479), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n671), .B2(new_n483), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n671), .A2(new_n264), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n453), .A2(new_n264), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n474), .A2(KEYINPUT38), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n400), .A2(new_n426), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n418), .B1(new_n472), .B2(new_n473), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n467), .A2(new_n468), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n690), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n481), .A2(new_n482), .B1(new_n432), .B2(new_n484), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n696), .A2(new_n697), .B1(new_n433), .B2(new_n440), .ZN(new_n698));
  INV_X1    g497(.A(new_n620), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n487), .A2(KEYINPUT44), .A3(new_n620), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  INV_X1    g502(.A(new_n543), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n540), .B1(new_n532), .B2(new_n534), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n542), .A2(KEYINPUT109), .A3(new_n543), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n644), .A3(new_n669), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n400), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n620), .A2(new_n544), .A3(new_n668), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT108), .Z(new_n713));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n644), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n549), .A3(new_n434), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(G1328gat));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n545), .A3(new_n675), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT46), .Z(new_n719));
  INV_X1    g518(.A(new_n675), .ZN(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n710), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1329gat));
  INV_X1    g521(.A(new_n483), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n700), .A2(new_n701), .A3(new_n723), .A4(new_n709), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT47), .B1(new_n725), .B2(KEYINPUT110), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n714), .A2(new_n552), .A3(new_n439), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n725), .B(new_n727), .C1(KEYINPUT110), .C2(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1330gat));
  NOR2_X1   g530(.A1(new_n264), .A2(new_n554), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n700), .A2(new_n701), .A3(new_n709), .A4(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n714), .A2(new_n484), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(G50gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n620), .A2(new_n544), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n644), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(KEYINPUT111), .A3(new_n669), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n668), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n487), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n487), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n400), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n489), .ZN(G1332gat));
  OAI22_X1  g549(.A1(new_n748), .A2(new_n720), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT49), .B(G64gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n745), .A2(new_n675), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1333gat));
  NAND3_X1  g553(.A1(new_n745), .A2(new_n747), .A3(new_n723), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G71gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n745), .A2(new_n747), .A3(new_n496), .A4(new_n439), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n748), .A2(new_n264), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n258), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n583), .A2(new_n585), .ZN(new_n764));
  INV_X1    g563(.A(new_n544), .ZN(new_n765));
  INV_X1    g564(.A(new_n644), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n668), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n702), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n770), .B2(new_n400), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n487), .A2(new_n620), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n768), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n698), .A2(new_n699), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n434), .A2(new_n583), .A3(new_n585), .A4(new_n669), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n771), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n720), .A2(G92gat), .A3(new_n668), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n700), .A2(new_n701), .A3(new_n675), .A4(new_n769), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(KEYINPUT114), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n775), .B2(new_n767), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n698), .A2(new_n772), .A3(new_n699), .A4(new_n768), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n781), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(G92gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n787), .A2(new_n793), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n770), .B2(new_n483), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n479), .A2(G99gat), .A3(new_n668), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n778), .B2(new_n796), .ZN(G1338gat));
  NOR3_X1   g596(.A1(new_n264), .A2(G106gat), .A3(new_n668), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n788), .B2(new_n789), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n700), .A2(new_n701), .A3(new_n484), .A4(new_n769), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n804), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n644), .A2(G113gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT119), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n656), .A2(new_n655), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT10), .B1(new_n650), .B2(KEYINPUT103), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n659), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n648), .B1(new_n657), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n810), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n657), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n649), .B1(new_n819), .B2(new_n815), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n665), .A2(new_n667), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n630), .B1(new_n629), .B2(new_n632), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n638), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n643), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n644), .A2(new_n824), .B1(new_n668), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n699), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n615), .B2(new_n619), .ZN(new_n831));
  INV_X1    g630(.A(new_n824), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n708), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n766), .A2(new_n620), .A3(new_n544), .A4(new_n669), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n809), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n372), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n737), .A2(new_n644), .A3(new_n668), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n829), .A2(new_n699), .B1(new_n831), .B2(new_n832), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(KEYINPUT116), .C1(new_n839), .C2(new_n708), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n837), .A3(new_n434), .A4(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT117), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(new_n720), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n842), .B2(new_n720), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n808), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n836), .A2(new_n840), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n400), .A3(new_n675), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n484), .A2(new_n479), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n644), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n851), .ZN(G1340gat));
  NOR2_X1   g651(.A1(new_n668), .A2(new_n322), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n844), .B2(new_n845), .ZN(new_n854));
  OAI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n668), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  NOR2_X1   g655(.A1(new_n544), .A2(G127gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n720), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n708), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1342gat));
  NOR2_X1   g660(.A1(new_n699), .A2(G134gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n720), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850), .B2(new_n699), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n842), .A2(new_n720), .A3(new_n862), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n863), .A2(new_n869), .A3(KEYINPUT56), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n864), .B(new_n865), .C1(new_n868), .C2(new_n870), .ZN(G1343gat));
  NAND3_X1  g670(.A1(new_n483), .A2(new_n434), .A3(new_n720), .ZN(new_n872));
  INV_X1    g671(.A(new_n839), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n835), .B1(new_n873), .B2(new_n544), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n874), .A2(new_n875), .A3(new_n264), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n836), .A2(new_n484), .A3(new_n840), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n875), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(KEYINPUT121), .A3(new_n875), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n872), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n206), .B1(new_n882), .B2(new_n766), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n723), .A2(new_n264), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n848), .A2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(G141gat), .A3(new_n644), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT58), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n886), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n644), .B(new_n872), .C1(new_n880), .C2(new_n881), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n206), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(G1344gat));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n208), .C1(new_n882), .C2(new_n669), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n894));
  NOR2_X1   g693(.A1(new_n873), .A2(KEYINPUT123), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n544), .B1(new_n839), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n838), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n875), .A3(new_n484), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n877), .A2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n901), .A2(new_n668), .A3(new_n872), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n669), .A2(new_n208), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n893), .A2(new_n903), .B1(new_n885), .B2(new_n904), .ZN(G1345gat));
  AND2_X1   g704(.A1(new_n882), .A2(new_n708), .ZN(new_n906));
  INV_X1    g705(.A(G155gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n765), .A2(new_n907), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n885), .B2(new_n908), .ZN(G1346gat));
  NOR2_X1   g708(.A1(new_n847), .A2(new_n400), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n675), .A2(new_n216), .A3(new_n699), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n884), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n882), .A2(new_n620), .ZN(new_n914));
  INV_X1    g713(.A(new_n216), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G1347gat));
  NAND2_X1  g715(.A1(new_n675), .A2(new_n400), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n847), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n849), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n644), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n847), .A2(new_n372), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n283), .A3(new_n766), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1348gat));
  OAI21_X1  g722(.A(G176gat), .B1(new_n919), .B2(new_n668), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n284), .A3(new_n669), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n919), .B2(new_n859), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n274), .A3(new_n765), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n275), .A3(new_n620), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n918), .A2(new_n849), .A3(new_n620), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(G190gat), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n932), .B2(G190gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  INV_X1    g736(.A(new_n877), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n723), .A2(new_n917), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n766), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n901), .A2(new_n723), .A3(new_n917), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n766), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  XOR2_X1   g748(.A(KEYINPUT126), .B(G204gat), .Z(new_n950));
  NAND2_X1  g749(.A1(new_n669), .A2(new_n950), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n940), .A2(new_n951), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n947), .A2(new_n669), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n954), .B(new_n955), .C1(new_n956), .C2(new_n950), .ZN(G1353gat));
  NAND4_X1  g756(.A1(new_n900), .A2(new_n899), .A3(new_n765), .A4(new_n939), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n544), .A2(G211gat), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n959), .A2(new_n960), .B1(new_n944), .B2(new_n961), .ZN(G1354gat));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n620), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G218gat), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n699), .A2(G218gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n944), .B2(new_n965), .ZN(G1355gat));
endmodule


