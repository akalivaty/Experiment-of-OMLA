//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT88), .B(G104), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n187), .B(new_n188), .Z(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  XNOR2_X1  g005(.A(G125), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT73), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(KEYINPUT16), .C1(new_n193), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n191), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n194), .B1(new_n193), .B2(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(KEYINPUT19), .B2(new_n192), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n203), .B2(new_n191), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G953), .ZN(new_n209));
  INV_X1    g023(.A(G237), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(new_n209), .A3(G214), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT86), .B(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(G953), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT86), .A2(G143), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(G214), .A3(new_n210), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n205), .B1(new_n217), .B2(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  AOI211_X1 g033(.A(KEYINPUT87), .B(new_n219), .C1(new_n213), .C2(new_n216), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n217), .A2(G131), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n204), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(G131), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n192), .A2(new_n191), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n201), .B2(new_n191), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n213), .B(new_n216), .C1(new_n225), .C2(new_n219), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n190), .B1(new_n223), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT89), .B1(new_n221), .B2(KEYINPUT17), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n236));
  NOR4_X1   g050(.A1(new_n218), .A2(new_n220), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  OAI221_X1 g052(.A(new_n236), .B1(G131), .B2(new_n217), .C1(new_n218), .C2(new_n220), .ZN(new_n239));
  INV_X1    g053(.A(new_n200), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n197), .A2(new_n191), .A3(new_n199), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n190), .B(new_n232), .C1(new_n238), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n224), .A2(KEYINPUT87), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n217), .A2(new_n205), .A3(G131), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT17), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n235), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n221), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n240), .A2(new_n241), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n222), .B1(new_n246), .B2(new_n247), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n236), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n231), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT90), .A3(new_n190), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n233), .B1(new_n245), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT20), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n257), .C2(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n245), .A2(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(new_n233), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT20), .B1(new_n259), .B2(KEYINPUT92), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n266), .B(new_n267), .C1(KEYINPUT92), .C2(new_n259), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n262), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n255), .A2(new_n190), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n245), .B2(new_n256), .ZN(new_n271));
  OAI21_X1  g085(.A(G475), .B1(new_n271), .B2(G902), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G116), .B(G122), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G128), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(new_n280), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n276), .B(new_n283), .C1(new_n286), .C2(new_n282), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n281), .B(new_n282), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n290));
  INV_X1    g104(.A(new_n274), .ZN(new_n291));
  OAI211_X1 g105(.A(G107), .B(new_n290), .C1(new_n291), .C2(KEYINPUT14), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n274), .A2(new_n275), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(KEYINPUT93), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n287), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n296), .B(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(G902), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n301), .B(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G952), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT94), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT94), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n206), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(G234), .B2(G237), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT21), .B(G898), .Z(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT95), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  AOI211_X1 g127(.A(new_n313), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT96), .B1(new_n273), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT96), .ZN(new_n319));
  INV_X1    g133(.A(new_n317), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n269), .A2(new_n319), .A3(new_n272), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n282), .B2(G137), .ZN(new_n324));
  INV_X1    g138(.A(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT11), .A3(G134), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n282), .A2(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n326), .A3(new_n219), .A4(new_n327), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n191), .A2(G143), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n279), .A2(G146), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT0), .A4(G128), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT0), .B(G128), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(KEYINPUT64), .A3(G131), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n332), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(KEYINPUT1), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G128), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n333), .B(new_n334), .C1(KEYINPUT1), .C2(new_n277), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n327), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n282), .A2(G137), .ZN(new_n348));
  OAI21_X1  g162(.A(G131), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n331), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n341), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT30), .ZN(new_n352));
  INV_X1    g166(.A(G119), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G116), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n289), .A2(G119), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT2), .B(G113), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n350), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT65), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n332), .A2(new_n339), .A3(new_n363), .A4(new_n340), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n352), .B(new_n360), .C1(new_n365), .C2(KEYINPUT30), .ZN(new_n366));
  INV_X1    g180(.A(new_n360), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n351), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n214), .A2(G210), .A3(new_n210), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT27), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT26), .B(G101), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT31), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n373), .A2(KEYINPUT31), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT67), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n377), .A3(KEYINPUT31), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n368), .B1(new_n365), .B2(new_n367), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n372), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n375), .A2(new_n376), .A3(new_n378), .A4(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G472), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n313), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT32), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT69), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT69), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n387), .A2(KEYINPUT32), .A3(new_n388), .A4(new_n313), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n372), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n366), .A2(new_n368), .A3(new_n385), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT29), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT70), .B1(new_n351), .B2(new_n367), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n367), .B2(new_n351), .ZN(new_n400));
  INV_X1    g214(.A(new_n351), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT70), .A3(new_n360), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n383), .B1(new_n403), .B2(new_n382), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n372), .A2(KEYINPUT29), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n313), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G472), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n392), .A2(new_n394), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n277), .A2(KEYINPUT23), .A3(G119), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n353), .A2(G128), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n353), .A2(G128), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(KEYINPUT23), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(G110), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT24), .B(G110), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n412), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n414), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n227), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT74), .B1(new_n422), .B2(new_n200), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n240), .A2(new_n424), .A3(new_n227), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT75), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT72), .B1(new_n417), .B2(new_n420), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(G110), .B2(new_n413), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n417), .A2(KEYINPUT72), .A3(new_n420), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n252), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n427), .B1(new_n426), .B2(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G137), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n437), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n427), .B(new_n439), .C1(new_n426), .C2(new_n431), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT76), .B(KEYINPUT25), .C1(new_n441), .C2(G902), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n443));
  INV_X1    g257(.A(new_n434), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n432), .A3(new_n439), .ZN(new_n445));
  INV_X1    g259(.A(new_n440), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n298), .B1(G234), .B2(new_n313), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n442), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(G902), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n438), .B2(new_n440), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n409), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n313), .ZN(new_n459));
  INV_X1    g273(.A(G104), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT3), .B1(new_n460), .B2(G107), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n275), .A3(G104), .ZN(new_n463));
  INV_X1    g277(.A(G101), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(G107), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n460), .A2(G107), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n275), .A2(G104), .ZN(new_n468));
  OAI21_X1  g282(.A(G101), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT79), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n472), .A2(KEYINPUT10), .A3(new_n346), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n346), .A2(new_n470), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G101), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n480), .A2(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT4), .A3(new_n466), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n339), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n332), .A2(new_n340), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n475), .A2(new_n478), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(G110), .B(G140), .Z(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT77), .ZN(new_n487));
  INV_X1    g301(.A(new_n214), .ZN(new_n488));
  INV_X1    g302(.A(G227), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n487), .B(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n344), .A2(new_n345), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n473), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n476), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n484), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT80), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(KEYINPUT80), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n495), .B2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(KEYINPUT80), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n475), .A2(new_n478), .A3(new_n483), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n496), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n485), .ZN(new_n506));
  INV_X1    g320(.A(new_n491), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n459), .B1(new_n509), .B2(new_n458), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n502), .A2(new_n485), .A3(new_n498), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n492), .A2(new_n505), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G469), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n457), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n338), .A2(G125), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n346), .B2(G125), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT83), .B(G224), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n206), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT84), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n526), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT5), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n531), .B(G113), .C1(KEYINPUT5), .C2(new_n354), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n358), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n472), .A3(new_n474), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n481), .A2(new_n360), .A3(new_n482), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n539), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n538), .A3(new_n536), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n529), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n523), .A2(new_n525), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n522), .B1(new_n546), .B2(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n473), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n538), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n533), .A2(new_n470), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n548), .A2(new_n543), .A3(new_n549), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n554), .A2(new_n313), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G210), .B1(G237), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n556), .B(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n518), .A2(new_n520), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n322), .A2(new_n455), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G101), .ZN(G3));
  AND2_X1   g377(.A1(new_n387), .A2(new_n313), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n388), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n389), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n451), .A2(new_n453), .A3(new_n517), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n302), .A2(new_n313), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n301), .B2(new_n302), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n300), .B(KEYINPUT33), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n573), .B2(new_n302), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n556), .A2(new_n557), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n545), .A2(new_n558), .A3(new_n555), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n519), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n315), .ZN(new_n580));
  AND4_X1   g394(.A1(KEYINPUT98), .A2(new_n273), .A3(new_n576), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n574), .B(KEYINPUT97), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n269), .B2(new_n272), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT98), .B1(new_n583), .B2(new_n580), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n569), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT99), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT100), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(KEYINPUT20), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n266), .A2(new_n590), .A3(new_n258), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT101), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n266), .A2(new_n593), .A3(new_n590), .A4(new_n258), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n262), .A3(new_n263), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n304), .ZN(new_n596));
  AND4_X1   g410(.A1(new_n272), .A2(new_n595), .A3(new_n596), .A4(new_n580), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n569), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NAND2_X1  g414(.A1(new_n426), .A2(new_n431), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n439), .A2(KEYINPUT36), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n452), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT102), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n451), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n567), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n322), .A2(new_n561), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT37), .B(G110), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G12));
  INV_X1    g425(.A(G900), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n309), .B1(new_n314), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND4_X1   g428(.A1(new_n272), .A2(new_n595), .A3(new_n596), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n392), .A2(new_n408), .A3(new_n394), .ZN(new_n616));
  INV_X1    g430(.A(new_n579), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n518), .B1(new_n451), .B2(new_n605), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  XNOR2_X1  g434(.A(new_n560), .B(KEYINPUT38), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n621), .A2(new_n304), .A3(new_n520), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n613), .B(KEYINPUT39), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n517), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT40), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n624), .A2(KEYINPUT40), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n607), .A2(new_n622), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n392), .A2(new_n394), .ZN(new_n628));
  INV_X1    g442(.A(new_n403), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n313), .B1(new_n629), .B2(new_n372), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n366), .A2(new_n368), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n372), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n395), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n627), .A2(new_n273), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(G143), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G45));
  AOI211_X1 g453(.A(new_n613), .B(new_n582), .C1(new_n269), .C2(new_n272), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n616), .A3(new_n617), .A4(new_n618), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G146), .ZN(G48));
  NAND2_X1  g456(.A1(new_n503), .A2(new_n508), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n313), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G469), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n509), .A2(new_n458), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n647));
  OR3_X1    g461(.A1(new_n509), .A2(KEYINPUT104), .A3(new_n458), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n456), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n409), .A2(new_n454), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n581), .B2(new_n584), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT41), .B(G113), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT105), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(G15));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n597), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G116), .ZN(G18));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n579), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n607), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n322), .A2(new_n616), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT106), .B(G119), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G21));
  NAND2_X1  g477(.A1(new_n404), .A2(new_n385), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n374), .A3(new_n376), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n388), .A3(new_n313), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n566), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n454), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n617), .A2(new_n596), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n649), .A2(new_n316), .A3(new_n456), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n669), .B(new_n670), .C1(new_n272), .C2(new_n269), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G122), .ZN(G24));
  NAND3_X1  g487(.A1(new_n273), .A2(new_n576), .A3(new_n614), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT107), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n583), .A2(new_n676), .A3(new_n614), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n566), .A2(new_n658), .A3(new_n606), .A4(new_n666), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G125), .ZN(G27));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n677), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n454), .B1(new_n408), .B2(new_n391), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n515), .A2(KEYINPUT108), .A3(G469), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n510), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT108), .B1(new_n515), .B2(G469), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n456), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n560), .A2(new_n519), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n454), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n616), .A2(new_n692), .A3(new_n688), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n675), .A3(new_n677), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G131), .ZN(G33));
  NAND2_X1  g514(.A1(new_n693), .A2(new_n615), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G134), .ZN(G36));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n704));
  INV_X1    g518(.A(new_n389), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n606), .B1(new_n565), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n269), .A2(new_n272), .A3(new_n576), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n269), .A2(KEYINPUT43), .A3(new_n272), .A4(new_n576), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n704), .B(new_n706), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n703), .B1(new_n711), .B2(new_n687), .ZN(new_n712));
  INV_X1    g526(.A(new_n687), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n710), .ZN(new_n714));
  INV_X1    g528(.A(new_n706), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(KEYINPUT110), .B(new_n713), .C1(new_n716), .C2(new_n704), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n458), .B1(new_n514), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT45), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n459), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n646), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n723), .B(new_n459), .C1(new_n719), .C2(new_n720), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n456), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n623), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n716), .B2(new_n704), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n712), .A2(new_n717), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G137), .ZN(G39));
  NAND2_X1  g544(.A1(new_n454), .A2(new_n713), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT47), .B(new_n456), .C1(new_n722), .C2(new_n724), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n409), .A3(new_n640), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G140), .ZN(G42));
  NAND4_X1  g551(.A1(new_n692), .A2(new_n621), .A3(new_n519), .A4(new_n456), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n649), .B(KEYINPUT49), .Z(new_n739));
  OR4_X1    g553(.A1(new_n636), .A2(new_n738), .A3(new_n707), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n669), .B1(new_n269), .B2(new_n272), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n606), .A2(new_n686), .A3(new_n613), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n636), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n679), .A2(new_n619), .A3(new_n641), .A4(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n273), .A2(new_n576), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n273), .B2(new_n304), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n560), .A2(new_n315), .A3(new_n520), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n567), .A2(new_n568), .A3(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n749), .A2(new_n751), .B1(new_n671), .B2(new_n668), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n562), .A3(new_n609), .A4(new_n661), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n652), .A2(new_n656), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n687), .A2(new_n596), .A3(new_n613), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n595), .A2(new_n755), .A3(new_n272), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT111), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n595), .A2(new_n755), .A3(new_n758), .A4(new_n272), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n616), .A3(new_n618), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n667), .A2(new_n607), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n688), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n701), .B(new_n760), .C1(new_n681), .C2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n753), .A2(new_n754), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n679), .A2(new_n619), .A3(new_n641), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n679), .A2(new_n619), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n744), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n747), .A2(new_n699), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT112), .ZN(new_n772));
  AND4_X1   g586(.A1(KEYINPUT53), .A2(new_n747), .A3(new_n699), .A4(new_n764), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n771), .B1(new_n773), .B2(KEYINPUT112), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n741), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n308), .ZN(new_n776));
  INV_X1    g590(.A(new_n636), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n650), .A2(new_n687), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n692), .A3(new_n309), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n714), .A2(new_n309), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n668), .ZN(new_n781));
  OAI221_X1 g595(.A(new_n776), .B1(new_n779), .B2(new_n748), .C1(new_n781), .C2(new_n659), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n778), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n682), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT48), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT48), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n650), .A2(KEYINPUT114), .A3(new_n519), .ZN(new_n789));
  OAI21_X1  g603(.A(KEYINPUT114), .B1(new_n650), .B2(new_n519), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n621), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT115), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT50), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n761), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n779), .A2(new_n273), .A3(new_n576), .ZN(new_n795));
  INV_X1    g609(.A(new_n781), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n733), .A2(new_n734), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n456), .B1(new_n649), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n798), .B2(new_n649), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n687), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n795), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n793), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT51), .A4(new_n802), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n788), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n769), .A2(KEYINPUT53), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n747), .A2(new_n770), .A3(new_n764), .A4(new_n699), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT54), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n775), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(G952), .A2(G953), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n740), .B1(new_n811), .B2(new_n812), .ZN(G75));
  NAND4_X1  g627(.A1(new_n808), .A2(G210), .A3(G902), .A4(new_n809), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n544), .A2(new_n541), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n530), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n815), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n214), .A2(G952), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n820), .A2(KEYINPUT117), .A3(new_n822), .A4(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(G51));
  XNOR2_X1  g643(.A(new_n459), .B(KEYINPUT57), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n808), .A2(new_n809), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n741), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(new_n810), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n643), .B(KEYINPUT118), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n831), .A2(new_n313), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n720), .A3(new_n719), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n823), .B1(new_n835), .B2(new_n837), .ZN(G54));
  NAND3_X1  g652(.A1(new_n836), .A2(KEYINPUT58), .A3(G475), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n257), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n824), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n839), .A2(new_n257), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(G60));
  XOR2_X1   g657(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n570), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n573), .B(new_n845), .C1(new_n832), .C2(new_n810), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n824), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n775), .B2(new_n810), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n572), .B2(new_n848), .ZN(G63));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n298), .A2(new_n313), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n808), .A2(new_n809), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n823), .B1(new_n853), .B2(new_n441), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n808), .A2(new_n603), .A3(new_n809), .A4(new_n852), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n854), .A2(new_n858), .A3(new_n859), .A4(new_n855), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(G66));
  OR2_X1    g677(.A1(new_n753), .A2(new_n754), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n214), .ZN(new_n865));
  INV_X1    g679(.A(new_n527), .ZN(new_n866));
  OAI21_X1  g680(.A(G953), .B1(new_n312), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n865), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT123), .ZN(new_n873));
  INV_X1    g687(.A(G898), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n817), .B1(new_n874), .B2(new_n488), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n873), .B(new_n875), .ZN(G69));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n488), .B1(new_n489), .B2(new_n612), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n766), .A2(new_n637), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT62), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n624), .A2(new_n687), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n749), .A2(new_n455), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(new_n736), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n766), .A2(new_n884), .A3(new_n637), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n883), .A3(new_n729), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n352), .B1(new_n365), .B2(KEYINPUT30), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n203), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n488), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n682), .A2(new_n623), .A3(new_n742), .A4(new_n726), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n701), .A2(new_n736), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n765), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n729), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n694), .A2(new_n696), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT109), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n690), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n214), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n214), .A2(G900), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n888), .B1(new_n904), .B2(KEYINPUT125), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n699), .A2(new_n729), .A3(new_n895), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n906), .B2(new_n214), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n892), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n877), .B(new_n878), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n878), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n910), .B2(new_n877), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n889), .B1(new_n907), .B2(new_n908), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT125), .B(new_n902), .C1(new_n906), .C2(new_n214), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n891), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n917), .B2(KEYINPUT124), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(G72));
  NAND2_X1  g734(.A1(G472), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT63), .Z(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n886), .B2(new_n864), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n633), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT127), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n632), .A2(new_n397), .A3(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n772), .B2(new_n774), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n906), .A2(new_n864), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n397), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n925), .A2(new_n927), .A3(new_n823), .A4(new_n929), .ZN(G57));
endmodule


