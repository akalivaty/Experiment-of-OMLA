//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT12), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n190), .A2(KEYINPUT11), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  AND4_X1   g008(.A1(KEYINPUT67), .A2(new_n193), .A3(new_n194), .A4(G134), .ZN(new_n195));
  AOI22_X1  g009(.A1(KEYINPUT67), .A2(new_n193), .B1(new_n194), .B2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(new_n192), .C1(new_n195), .C2(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(G107), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(new_n207), .C1(new_n208), .C2(new_n203), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT84), .B(G101), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n212));
  INV_X1    g026(.A(new_n207), .ZN(new_n213));
  OAI21_X1  g027(.A(G101), .B1(new_n213), .B2(new_n208), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G143), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n219), .B2(G143), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(KEYINPUT65), .A3(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n220), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n220), .B1(new_n216), .B2(new_n217), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT70), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n224), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n214), .B1(new_n209), .B2(new_n210), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT85), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n215), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n240), .A2(KEYINPUT86), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n218), .A2(new_n223), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n221), .A2(G146), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(G128), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n220), .A2(new_n222), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n238), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n240), .B2(KEYINPUT86), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n189), .B(new_n202), .C1(new_n241), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n241), .A2(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT12), .A3(new_n201), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT87), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT12), .B1(new_n253), .B2(new_n201), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n215), .A2(new_n239), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n229), .A2(new_n236), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n242), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(KEYINPUT10), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n209), .A2(G101), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT0), .A4(G128), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n243), .B1(new_n226), .B2(new_n227), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n263), .A2(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n248), .A2(KEYINPUT10), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n262), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n202), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n258), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n273), .A2(new_n202), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n274), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n187), .B(new_n188), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n258), .A2(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(KEYINPUT88), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT88), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n290), .A3(new_n283), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(G469), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(G469), .A2(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  OAI21_X1  g109(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n237), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n268), .A2(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(KEYINPUT91), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(KEYINPUT91), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G953), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G224), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT90), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n306), .B(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT2), .B(G113), .Z(new_n312));
  XNOR2_X1  g126(.A(G116), .B(G119), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n270), .A3(new_n264), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n316), .A2(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(KEYINPUT5), .ZN(new_n322));
  INV_X1    g136(.A(G116), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n322), .B(G113), .C1(KEYINPUT5), .C2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n259), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G122), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT89), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n328), .A2(KEYINPUT6), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n327), .A3(new_n329), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(KEYINPUT6), .B1(new_n328), .B2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n311), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n309), .A2(KEYINPUT7), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n303), .B(new_n335), .Z(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n321), .A2(new_n326), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n238), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n327), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n329), .B(KEYINPUT8), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G902), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G210), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n334), .A2(new_n345), .A3(new_n343), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n299), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G122), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G116), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n323), .A2(G122), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT95), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(KEYINPUT95), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n204), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n354), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n355), .B(KEYINPUT14), .ZN(new_n362));
  OAI21_X1  g176(.A(G107), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n221), .A2(G128), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT96), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT70), .B(G128), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G134), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n191), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n360), .A2(KEYINPUT98), .A3(new_n363), .A4(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n354), .A2(new_n355), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G107), .B1(new_n376), .B2(new_n357), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n371), .A2(new_n363), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n365), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n367), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n365), .A2(new_n381), .ZN(new_n384));
  OAI21_X1  g198(.A(G134), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n370), .B(KEYINPUT97), .Z(new_n386));
  NOR3_X1   g200(.A1(new_n358), .A2(new_n204), .A3(new_n359), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n377), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n295), .A2(new_n390), .A3(G953), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT99), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n380), .A2(new_n388), .A3(new_n392), .ZN(new_n395));
  AOI21_X1  g209(.A(G902), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n396), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(G237), .A2(G953), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G214), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(G143), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT92), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  XNOR2_X1  g222(.A(G125), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n219), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n300), .A2(KEYINPUT77), .A3(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n410), .B1(new_n414), .B2(new_n219), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n408), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n404), .B(G131), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n300), .A2(KEYINPUT16), .A3(G140), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT78), .Z(new_n421));
  INV_X1    g235(.A(new_n414), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT16), .ZN(new_n423));
  OAI211_X1 g237(.A(G146), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n219), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n404), .A2(new_n418), .A3(new_n199), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n419), .A2(new_n424), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n416), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n206), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n424), .B(KEYINPUT79), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n409), .A2(KEYINPUT19), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n414), .B2(KEYINPUT19), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G146), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n417), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n416), .B(new_n433), .C1(new_n434), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT20), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n432), .A2(new_n444), .A3(new_n439), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n433), .A2(KEYINPUT93), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n429), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n429), .A2(new_n446), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n188), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n443), .A2(new_n445), .B1(new_n449), .B2(G475), .ZN(new_n450));
  NAND2_X1  g264(.A1(G234), .A2(G237), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(G952), .A3(new_n307), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(G902), .A3(G953), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT100), .Z(new_n457));
  NAND3_X1  g271(.A1(new_n401), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n297), .A2(new_n350), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n201), .A2(new_n269), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n191), .A2(G137), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n194), .A2(G134), .ZN(new_n463));
  OAI21_X1  g277(.A(G131), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n261), .A2(new_n200), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n319), .B1(new_n466), .B2(KEYINPUT74), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(KEYINPUT74), .B2(new_n466), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n200), .A2(new_n464), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n471), .A2(KEYINPUT68), .B1(new_n260), .B2(new_n242), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n198), .A2(new_n200), .B1(new_n268), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n472), .A2(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(new_n318), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n319), .A2(new_n466), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n402), .A2(G210), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G101), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n461), .A2(new_n465), .A3(KEYINPUT30), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n319), .B(new_n490), .C1(new_n477), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n479), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n486), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT73), .A4(new_n486), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n489), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n495), .A2(new_n489), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n488), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G472), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n488), .B(KEYINPUT75), .C1(new_n499), .C2(new_n500), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n188), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT32), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n504), .A4(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n493), .A2(new_n494), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n512), .A2(new_n486), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n514), .C1(new_n481), .C2(new_n487), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n466), .B(new_n318), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n469), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n469), .B2(new_n468), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n487), .A2(new_n514), .ZN(new_n519));
  AOI21_X1  g333(.A(G902), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n504), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n366), .A2(G119), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(G119), .B2(new_n231), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT24), .B(G110), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n528));
  NOR2_X1   g342(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n529));
  INV_X1    g343(.A(G119), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n528), .A2(new_n529), .B1(new_n530), .B2(G128), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT23), .ZN(new_n532));
  OAI221_X1 g346(.A(new_n531), .B1(G119), .B2(new_n231), .C1(new_n524), .C2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n527), .B1(new_n533), .B2(G110), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n410), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n434), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n426), .A2(new_n424), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(G110), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n525), .C2(new_n526), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT22), .B(G137), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n307), .A2(G221), .A3(G234), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n536), .A2(new_n539), .A3(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT82), .ZN(new_n548));
  INV_X1    g362(.A(G234), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n549), .B2(G217), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT25), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n546), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G217), .B1(new_n549), .B2(G902), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n460), .B1(new_n523), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n521), .B1(new_n507), .B2(new_n510), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(KEYINPUT83), .A3(new_n561), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n459), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n210), .ZN(G3));
  NAND3_X1  g381(.A1(new_n503), .A2(new_n188), .A3(new_n505), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n506), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n294), .A2(new_n296), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n562), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n349), .A2(new_n457), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n396), .A2(G478), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n394), .A2(new_n395), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT33), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n397), .A2(G902), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n576), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n450), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT34), .B(G104), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  NAND3_X1  g404(.A1(new_n400), .A2(new_n450), .A3(new_n457), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT102), .Z(new_n592));
  NOR2_X1   g406(.A1(new_n297), .A2(new_n350), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n571), .A4(new_n562), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT35), .B(G107), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT103), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n594), .B(new_n596), .ZN(G9));
  INV_X1    g411(.A(new_n459), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n540), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n550), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n560), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n570), .A2(KEYINPUT104), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT104), .B1(new_n570), .B2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT37), .B(G110), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G12));
  NAND4_X1  g423(.A1(new_n294), .A2(new_n349), .A3(new_n296), .A4(new_n602), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n564), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n450), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n401), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n455), .A2(G900), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n452), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  XNOR2_X1  g433(.A(new_n615), .B(KEYINPUT39), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n572), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT40), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n625), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n497), .A2(new_n498), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n516), .A2(new_n486), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n188), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n511), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n347), .A2(new_n348), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n635), .B(KEYINPUT38), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n400), .A2(new_n612), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n636), .A2(new_n299), .A3(new_n602), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n626), .A2(new_n629), .A3(new_n634), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G143), .ZN(G45));
  INV_X1    g454(.A(new_n615), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n585), .A2(new_n450), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n611), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  NOR2_X1   g458(.A1(new_n282), .A2(new_n284), .ZN(new_n645));
  OAI21_X1  g459(.A(G469), .B1(new_n645), .B2(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n285), .A3(new_n296), .ZN(new_n647));
  NOR4_X1   g461(.A1(new_n564), .A2(new_n587), .A3(new_n561), .A4(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT41), .B(G113), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G15));
  NOR2_X1   g464(.A1(new_n564), .A2(new_n561), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n647), .A2(new_n350), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n651), .A2(new_n592), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n323), .ZN(G18));
  NOR3_X1   g468(.A1(new_n647), .A2(new_n350), .A3(new_n603), .ZN(new_n655));
  INV_X1    g469(.A(new_n458), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n564), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n530), .ZN(G21));
  NOR3_X1   g473(.A1(new_n647), .A2(new_n574), .A3(new_n637), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n518), .A2(KEYINPUT106), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n518), .A2(KEYINPUT106), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n661), .A2(new_n662), .A3(new_n486), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n499), .A2(new_n500), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n504), .B(new_n188), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n569), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n562), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  NAND3_X1  g482(.A1(new_n655), .A2(new_n642), .A3(new_n666), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G125), .ZN(G27));
  NOR2_X1   g484(.A1(new_n635), .A2(new_n299), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n297), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n651), .A2(new_n642), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT42), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G131), .ZN(G33));
  XOR2_X1   g490(.A(new_n616), .B(KEYINPUT107), .Z(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n651), .A3(new_n673), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G134), .ZN(G36));
  INV_X1    g493(.A(new_n285), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n287), .A2(new_n291), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(KEYINPUT45), .ZN(new_n682));
  OAI21_X1  g496(.A(G469), .B1(new_n681), .B2(KEYINPUT45), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n293), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n296), .A3(new_n620), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n583), .A2(new_n584), .ZN(new_n689));
  INV_X1    g503(.A(new_n576), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n450), .B(KEYINPUT109), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n585), .A2(new_n612), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n693), .B(KEYINPUT43), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n694), .B2(KEYINPUT108), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n570), .A3(new_n602), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n672), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n688), .B(new_n701), .C1(new_n700), .C2(new_n699), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G137), .ZN(G39));
  NAND2_X1  g517(.A1(new_n687), .A2(new_n296), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n687), .A2(KEYINPUT47), .A3(new_n296), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n564), .A2(new_n561), .A3(new_n642), .A4(new_n671), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT110), .B(G140), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G42));
  INV_X1    g526(.A(new_n588), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n566), .A2(new_n713), .A3(KEYINPUT112), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n523), .A2(new_n460), .A3(new_n562), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT83), .B1(new_n564), .B2(new_n561), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n598), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n715), .B1(new_n718), .B2(new_n588), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n400), .B(KEYINPUT113), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n612), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n575), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n573), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n605), .B2(new_n606), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n714), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n714), .A2(new_n719), .A3(KEYINPUT114), .A4(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n667), .B1(new_n564), .B2(new_n657), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n648), .A3(new_n653), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n675), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n350), .A2(new_n637), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n602), .A2(new_n641), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n634), .A2(new_n572), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n618), .A2(new_n643), .A3(new_n669), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n666), .A2(new_n642), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n741), .A2(new_n655), .B1(new_n611), .B2(new_n617), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT52), .A3(new_n643), .A4(new_n736), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n720), .A2(new_n450), .A3(new_n615), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n740), .B1(new_n564), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n602), .A3(new_n673), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n678), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AND4_X1   g564(.A1(KEYINPUT53), .A2(new_n729), .A3(new_n733), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n727), .B2(new_n728), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT53), .B1(new_n752), .B2(new_n733), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT54), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n732), .A2(KEYINPUT115), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n732), .B2(KEYINPUT115), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n732), .B(new_n749), .C1(new_n727), .C2(new_n728), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(KEYINPUT53), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n762));
  INV_X1    g576(.A(new_n452), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n696), .A2(new_n763), .A3(new_n698), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n666), .A2(new_n562), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n647), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n636), .A2(new_n299), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(KEYINPUT50), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n768), .A3(new_n765), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n671), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n774), .A2(new_n634), .A3(new_n452), .A4(new_n561), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n450), .A3(new_n585), .ZN(new_n776));
  INV_X1    g590(.A(new_n774), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n764), .A2(new_n602), .A3(new_n666), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n296), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n646), .A2(new_n285), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n706), .A2(new_n707), .A3(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n671), .A3(new_n766), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n779), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n762), .B(new_n781), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n786), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n671), .A3(new_n766), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n788), .B(new_n789), .C1(new_n780), .C2(KEYINPUT51), .ZN(new_n790));
  INV_X1    g604(.A(G952), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n791), .B(G953), .C1(new_n766), .C2(new_n652), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n764), .A2(new_n651), .A3(new_n777), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT48), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n775), .A2(new_n586), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n787), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n754), .A2(new_n761), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(new_n307), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n693), .A2(new_n299), .A3(new_n561), .A4(new_n782), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n636), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n646), .A2(new_n285), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT49), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n802), .A2(new_n634), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n800), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(G75));
  AND3_X1   g626(.A1(new_n752), .A2(new_n755), .A3(new_n757), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n753), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n188), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(KEYINPUT119), .A3(G210), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n752), .A2(new_n733), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n756), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n758), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(G210), .A3(G902), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n333), .A2(new_n331), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n311), .ZN(new_n824));
  XOR2_X1   g638(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n816), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n307), .A2(G952), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT121), .Z(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n820), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n832), .B1(new_n834), .B2(new_n826), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n829), .A2(new_n835), .ZN(G51));
  INV_X1    g650(.A(new_n761), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n759), .B1(new_n818), .B2(new_n758), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n293), .B(KEYINPUT57), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n839), .A2(new_n840), .B1(new_n284), .B2(new_n282), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n682), .A2(new_n683), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT122), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n815), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n830), .B1(new_n841), .B2(new_n844), .ZN(G54));
  NAND2_X1  g659(.A1(KEYINPUT58), .A2(G475), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT123), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n815), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n440), .ZN(new_n849));
  INV_X1    g663(.A(new_n830), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n848), .B2(new_n440), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(G60));
  NAND2_X1  g666(.A1(G478), .A2(G902), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT59), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n583), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n831), .B1(new_n839), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n754), .A2(new_n761), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n583), .B1(new_n857), .B2(new_n854), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(G63));
  INV_X1    g673(.A(new_n548), .ZN(new_n860));
  NAND2_X1  g674(.A1(G217), .A2(G902), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT60), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n814), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n819), .A2(new_n600), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n831), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(G66));
  AOI21_X1  g682(.A(new_n307), .B1(new_n454), .B2(G224), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n729), .A2(new_n731), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n307), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n823), .B1(G898), .B2(new_n307), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n871), .B(new_n872), .Z(G69));
  INV_X1    g687(.A(new_n710), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n688), .A2(new_n651), .A3(new_n734), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n702), .A2(new_n678), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n742), .A2(new_n643), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n675), .A4(new_n877), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(G953), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n490), .B1(new_n477), .B2(new_n492), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(new_n436), .Z(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(G900), .B2(G953), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n639), .A2(new_n877), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n671), .B1(new_n721), .B2(new_n586), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n624), .A2(new_n625), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n563), .B2(new_n565), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n887), .A2(new_n702), .A3(new_n874), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n307), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n882), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n880), .B1(new_n879), .B2(new_n883), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n884), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(G900), .ZN(new_n897));
  OAI21_X1  g711(.A(G953), .B1(new_n276), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT124), .Z(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n879), .B2(new_n883), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n901), .A2(KEYINPUT125), .A3(new_n893), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT125), .B1(new_n901), .B2(new_n893), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n896), .A2(new_n898), .B1(new_n902), .B2(new_n903), .ZN(G72));
  NOR2_X1   g718(.A1(new_n751), .A2(new_n753), .ZN(new_n905));
  NAND2_X1  g719(.A1(G472), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT63), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n630), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n513), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT127), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n878), .B2(new_n870), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n487), .A3(new_n512), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n850), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n907), .B1(new_n891), .B2(new_n870), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n512), .A2(new_n487), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n912), .B(new_n915), .C1(new_n916), .C2(new_n917), .ZN(G57));
endmodule


