//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(G1gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G22gat), .Z(new_n206));
  OR2_X1    g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n202), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT89), .A3(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n209), .B(G8gat), .C1(KEYINPUT89), .C2(new_n208), .ZN(new_n210));
  AOI21_X1  g009(.A(G8gat), .B1(new_n207), .B2(KEYINPUT90), .ZN(new_n211));
  OR3_X1    g010(.A1(new_n205), .A2(KEYINPUT90), .A3(new_n206), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n224), .A2(new_n216), .A3(new_n215), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n214), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n210), .A2(new_n213), .B1(new_n226), .B2(new_n225), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n210), .A2(new_n213), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(new_n227), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT18), .A4(new_n232), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  INV_X1    g042(.A(G197gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT11), .B(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n235), .A2(new_n240), .A3(new_n248), .A4(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G8gat), .B(G36gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(G64gat), .B(G92gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n257), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G226gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G169gat), .ZN(new_n271));
  INV_X1    g070(.A(G176gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n274), .B(new_n275), .C1(new_n278), .C2(KEYINPUT26), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT27), .B(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT27), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT28), .B1(new_n286), .B2(KEYINPUT67), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n287), .B(new_n281), .C1(KEYINPUT67), .C2(new_n280), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n279), .A2(new_n283), .A3(new_n284), .A4(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n277), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT23), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n281), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  OAI221_X1 g095(.A(new_n293), .B1(new_n294), .B2(new_n295), .C1(new_n296), .C2(KEYINPUT66), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n275), .B1(new_n276), .B2(KEYINPUT23), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT25), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n293), .B1(new_n302), .B2(KEYINPUT64), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(KEYINPUT64), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT25), .B1(new_n276), .B2(KEYINPUT23), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n299), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n301), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n270), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n270), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n267), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n314), .ZN(new_n316));
  INV_X1    g115(.A(new_n267), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n316), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n256), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n267), .A3(new_n314), .ZN(new_n320));
  INV_X1    g119(.A(new_n256), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n316), .B2(new_n312), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(KEYINPUT30), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT30), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .A4(new_n321), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G141gat), .B(G148gat), .Z(new_n334));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT2), .ZN(new_n336));
  INV_X1    g135(.A(G155gat), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n335), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n334), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n335), .B(new_n339), .C1(new_n342), .C2(KEYINPUT2), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  INV_X1    g147(.A(G127gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT69), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(G113gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G120gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT1), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n347), .A2(G127gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n351), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT68), .ZN(new_n362));
  OR3_X1    g161(.A1(new_n347), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n362), .B(new_n363), .C1(KEYINPUT1), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n361), .A2(new_n365), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n341), .A2(new_n343), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n369), .A2(KEYINPUT75), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n361), .A2(new_n365), .A3(new_n343), .A4(new_n341), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n372), .A2(new_n375), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n368), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT39), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n333), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n367), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n344), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(new_n374), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n382), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n386), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT39), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n385), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT40), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n327), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT5), .B1(new_n392), .B2(new_n382), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g200(.A(new_n376), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n374), .A2(KEYINPUT4), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n367), .B(new_n382), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT73), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n405), .B(KEYINPUT5), .C1(new_n392), .C2(new_n382), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n368), .A2(new_n389), .ZN(new_n409));
  AND4_X1   g208(.A1(KEYINPUT77), .A2(new_n387), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT5), .B1(new_n378), .B2(new_n380), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT77), .B1(new_n411), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n409), .A3(new_n408), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(KEYINPUT86), .A3(new_n407), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n332), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n399), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT84), .B(new_n385), .C1(new_n394), .C2(new_n396), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n332), .B1(new_n390), .B2(KEYINPUT39), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n393), .B1(new_n381), .B2(new_n382), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n396), .B1(new_n427), .B2(KEYINPUT83), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n429), .A3(new_n398), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT85), .A4(new_n398), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n407), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n418), .B2(new_n419), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n437));
  AOI211_X1 g236(.A(new_n414), .B(new_n435), .C1(new_n418), .C2(new_n419), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n333), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n332), .B(new_n407), .C1(new_n410), .C2(new_n412), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n413), .A2(new_n333), .A3(new_n441), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n413), .A2(KEYINPUT87), .A3(new_n333), .A4(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT38), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n320), .A2(KEYINPUT37), .A3(new_n322), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT37), .B1(new_n320), .B2(new_n322), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n450), .B1(new_n453), .B2(new_n256), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n450), .B(new_n256), .C1(new_n451), .C2(new_n452), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n323), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n445), .A2(new_n448), .A3(new_n449), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G78gat), .B(G106gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT31), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT79), .B(G50gat), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n267), .B1(new_n463), .B2(new_n311), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n265), .B2(new_n266), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n344), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n468), .A2(KEYINPUT80), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n266), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n263), .B1(new_n261), .B2(new_n257), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n311), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n371), .B1(new_n474), .B2(new_n345), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT80), .B(new_n468), .C1(new_n475), .C2(new_n464), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n476), .A3(G22gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(G22gat), .B1(new_n471), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n462), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n476), .ZN(new_n481));
  INV_X1    g280(.A(G22gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(new_n485), .A3(new_n489), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n434), .A2(new_n458), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G227gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n269), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n310), .A2(new_n366), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n303), .B1(KEYINPUT64), .B2(new_n302), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n298), .B1(new_n496), .B2(new_n305), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n497), .A2(new_n308), .B1(new_n300), .B2(KEYINPUT25), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n369), .B1(new_n498), .B2(new_n289), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT33), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n494), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n310), .A2(new_n366), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n369), .A3(new_n289), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G43gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G71gat), .ZN(new_n510));
  INV_X1    g309(.A(G99gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n502), .A2(new_n508), .A3(KEYINPUT70), .A4(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT70), .B(new_n512), .C1(new_n506), .C2(KEYINPUT33), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n500), .A2(KEYINPUT32), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n505), .A3(new_n503), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n517), .A2(new_n519), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n513), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n513), .B2(new_n516), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT36), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT71), .ZN(new_n526));
  INV_X1    g325(.A(new_n516), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n514), .A2(new_n515), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n516), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(KEYINPUT36), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n324), .A2(new_n326), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n332), .B1(new_n420), .B2(new_n407), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n443), .A2(new_n536), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n436), .A2(new_n332), .A3(new_n442), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n491), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n492), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n523), .A2(new_n524), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n543), .A2(new_n535), .A3(new_n491), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n415), .A2(new_n421), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n443), .B1(new_n546), .B2(new_n333), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n448), .A2(new_n449), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n544), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n529), .A2(new_n532), .B1(new_n488), .B2(new_n490), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n535), .B(new_n550), .C1(new_n537), .C2(new_n538), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n253), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT20), .Z(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(KEYINPUT21), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n214), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n567));
  INV_X1    g366(.A(new_n565), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n563), .B1(new_n236), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n567), .B1(new_n566), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n556), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT94), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT19), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n566), .A2(new_n569), .ZN(new_n579));
  INV_X1    g378(.A(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n556), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n570), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n578), .B1(new_n573), .B2(new_n583), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT97), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n596), .A3(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n559), .B(new_n560), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n598), .A2(new_n561), .A3(new_n605), .A4(new_n599), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n598), .A2(new_n561), .A3(KEYINPUT10), .A4(new_n599), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n603), .A2(new_n606), .ZN(new_n615));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n228), .A2(new_n600), .ZN(new_n627));
  NAND3_X1  g426(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n598), .A2(new_n227), .A3(new_n599), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n627), .A2(new_n632), .A3(new_n628), .A4(new_n629), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n630), .A2(KEYINPUT98), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n635), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n587), .A2(new_n626), .A3(new_n644), .A4(KEYINPUT102), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n585), .A2(new_n586), .B1(new_n642), .B2(new_n641), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n647), .B2(new_n625), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n554), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n537), .A2(new_n538), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(KEYINPUT103), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n202), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n650), .A2(new_n535), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT16), .B(G8gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT105), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(KEYINPUT42), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n650), .B2(new_n535), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n662), .B1(new_n666), .B2(G8gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n659), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n667), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n650), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n670), .B2(new_n543), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n534), .A2(G15gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT106), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n670), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n650), .A2(new_n491), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  AOI21_X1  g476(.A(new_n644), .B1(new_n542), .B2(new_n553), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n587), .A2(new_n625), .A3(new_n253), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n652), .A2(new_n653), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n220), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n553), .A2(KEYINPUT108), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n549), .A2(new_n552), .A3(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n688), .A2(new_n690), .B1(new_n541), .B2(new_n492), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n687), .B1(new_n691), .B2(new_n644), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n680), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n654), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n686), .A2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n682), .A2(new_n221), .A3(new_n327), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n694), .B2(new_n535), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  INV_X1    g499(.A(new_n534), .ZN(new_n701));
  OAI21_X1  g500(.A(G43gat), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  INV_X1    g502(.A(G43gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n682), .A2(new_n704), .A3(new_n543), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n692), .A2(new_n540), .A3(new_n693), .A4(new_n680), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(G50gat), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n491), .A2(G50gat), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n679), .A2(new_n681), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI221_X4 g515(.A(new_n713), .B1(new_n709), .B2(KEYINPUT48), .C1(new_n710), .C2(G50gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  AOI21_X1  g517(.A(new_n689), .B1(new_n549), .B2(new_n552), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n549), .A2(new_n552), .A3(new_n689), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n542), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n647), .A2(new_n252), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n721), .A2(new_n625), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n683), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n327), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT49), .B(G64gat), .Z(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(G1333gat));
  NAND4_X1  g528(.A1(new_n721), .A2(new_n625), .A3(new_n534), .A4(new_n722), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(G71gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n721), .A2(new_n625), .A3(new_n722), .ZN(new_n732));
  INV_X1    g531(.A(new_n543), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n732), .A2(G71gat), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT110), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(G71gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n723), .A2(new_n736), .A3(new_n543), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n730), .A2(G71gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n735), .A2(KEYINPUT50), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT50), .B1(new_n735), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(G1334gat));
  NOR2_X1   g542(.A1(new_n732), .A2(new_n491), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT111), .B(G78gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n587), .A2(new_n252), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n692), .A2(new_n625), .A3(new_n693), .A4(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n589), .A3(new_n654), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n721), .A2(new_n643), .A3(new_n747), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n643), .A4(new_n747), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n626), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n683), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n749), .B1(new_n589), .B2(new_n755), .ZN(G1336gat));
  OAI21_X1  g555(.A(G92gat), .B1(new_n748), .B2(new_n535), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n625), .A2(new_n590), .A3(new_n327), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT112), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n757), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1337gat));
  NOR3_X1   g565(.A1(new_n748), .A2(new_n511), .A3(new_n701), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n754), .A2(new_n543), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n511), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  AOI21_X1  g569(.A(G106gat), .B1(new_n754), .B2(new_n540), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n540), .A2(G106gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n748), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n748), .A2(new_n772), .ZN(new_n775));
  AOI211_X1 g574(.A(new_n626), .B(new_n491), .C1(new_n752), .C2(new_n753), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n775), .B(KEYINPUT53), .C1(new_n776), .C2(G106gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1339gat));
  NOR3_X1   g577(.A1(new_n647), .A2(new_n625), .A3(new_n252), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n607), .A2(new_n611), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n780), .A2(KEYINPUT113), .A3(new_n616), .A4(new_n610), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n612), .B2(new_n613), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n612), .A2(new_n613), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n781), .B(KEYINPUT54), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n614), .A2(KEYINPUT54), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n624), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n614), .A2(new_n617), .A3(new_n624), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT55), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n232), .B1(new_n229), .B2(new_n231), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n236), .A2(new_n227), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(new_n230), .A3(new_n239), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n793), .B(new_n247), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n251), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n230), .B1(new_n214), .B2(new_n228), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n237), .A2(new_n239), .B1(new_n799), .B2(new_n232), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n793), .B1(new_n800), .B2(new_n247), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n587), .B1(new_n803), .B2(new_n643), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n790), .A2(new_n252), .A3(new_n791), .A4(new_n792), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n643), .B1(new_n625), .B2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n779), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n550), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n654), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n535), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n354), .A3(new_n252), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n803), .A2(new_n643), .ZN(new_n813));
  INV_X1    g612(.A(new_n587), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n807), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n779), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n683), .A3(new_n544), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n253), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n819), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n818), .B2(new_n626), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n625), .A2(new_n352), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT116), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n811), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1341gat));
  NOR3_X1   g625(.A1(new_n818), .A2(new_n349), .A3(new_n814), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n587), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT117), .Z(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n829), .B2(new_n349), .ZN(G1342gat));
  NAND2_X1  g629(.A1(new_n643), .A2(new_n535), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT118), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n347), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n818), .B2(new_n644), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n808), .A2(new_n491), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n654), .A2(new_n327), .A3(new_n534), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(G141gat), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(new_n844), .A3(new_n252), .ZN(new_n845));
  INV_X1    g644(.A(new_n842), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n808), .B2(new_n491), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n540), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n817), .B2(new_n540), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n808), .A2(new_n847), .A3(new_n491), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT120), .B(new_n842), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n252), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n845), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n844), .B1(new_n850), .B2(new_n252), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n845), .A2(KEYINPUT58), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n857), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(G1344gat));
  AOI22_X1  g660(.A1(new_n649), .A2(new_n253), .B1(new_n804), .B2(new_n807), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n847), .B1(new_n862), .B2(new_n491), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n626), .B1(new_n863), .B2(new_n849), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(KEYINPUT59), .A3(new_n842), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n626), .B1(new_n868), .B2(new_n854), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(KEYINPUT59), .ZN(new_n870));
  AOI21_X1  g669(.A(G148gat), .B1(new_n843), .B2(new_n625), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n870), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n871), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n843), .A2(new_n337), .A3(new_n587), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n814), .B1(new_n868), .B2(new_n854), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n337), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT121), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n873), .C1(new_n874), .C2(new_n337), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n654), .A2(G162gat), .A3(new_n534), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n841), .A2(new_n832), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n644), .B1(new_n868), .B2(new_n854), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n338), .ZN(G1347gat));
  NAND3_X1  g683(.A1(new_n817), .A2(new_n654), .A3(new_n327), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n809), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n271), .A3(new_n252), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n885), .A2(new_n540), .A3(new_n733), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n252), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n271), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n886), .B2(new_n625), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n626), .A2(new_n272), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n886), .A2(new_n587), .A3(new_n280), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n888), .A2(new_n587), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n285), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(G1350gat));
  AOI21_X1  g697(.A(new_n281), .B1(new_n888), .B2(new_n643), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT61), .Z(new_n900));
  NAND3_X1  g699(.A1(new_n886), .A2(new_n281), .A3(new_n643), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1351gat));
  NAND3_X1  g701(.A1(new_n654), .A2(new_n327), .A3(new_n701), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n808), .A3(new_n491), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n244), .A3(new_n252), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n253), .B(new_n903), .C1(new_n863), .C2(new_n849), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n244), .B2(new_n908), .ZN(G1352gat));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n625), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n903), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n864), .B2(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n913), .A2(new_n915), .A3(KEYINPUT126), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT126), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1353gat));
  NAND3_X1  g717(.A1(new_n906), .A2(new_n259), .A3(new_n587), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n863), .A2(new_n849), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n587), .A3(new_n914), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  AOI21_X1  g723(.A(G218gat), .B1(new_n906), .B2(new_n643), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n644), .A2(new_n260), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n914), .A3(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n925), .A2(KEYINPUT127), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT127), .B1(new_n925), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


