//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT69), .Z(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT71), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT71), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n478), .A2(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT72), .Z(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n472), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(new_n470), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n470), .A3(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n481), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n470), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n469), .A2(new_n472), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  AND3_X1   g086(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT74), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n521), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT75), .B1(new_n529), .B2(new_n518), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(G166));
  XOR2_X1   g106(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n516), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n509), .A2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT76), .B(G51), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  AOI22_X1  g117(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n521), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT78), .B(G52), .Z(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n510), .A2(new_n545), .B1(new_n516), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n521), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n510), .A2(new_n551), .B1(new_n516), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n521), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n535), .A2(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G166), .ZN(G303));
  OAI21_X1  g142(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n526), .A2(G87), .A3(new_n509), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NOR2_X1   g146(.A1(new_n512), .A2(new_n513), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n526), .A2(G86), .A3(new_n509), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G60), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n572), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n521), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n584), .B2(new_n583), .ZN(new_n586));
  AOI22_X1  g161(.A1(G47), .A2(new_n538), .B1(new_n535), .B2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n535), .A2(G92), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n572), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n538), .B2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n598), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g185(.A(KEYINPUT3), .B(G2104), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n474), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n490), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n492), .A2(G123), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n621), .ZN(G156));
  INV_X1    g197(.A(KEYINPUT14), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n626), .B2(new_n625), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n628), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n636), .A3(G14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT80), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT82), .B(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n640), .A2(new_n641), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n646), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n658), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n662), .C1(new_n655), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(G229));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NOR2_X1   g251(.A1(G303), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G16), .A2(G22), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n677), .A2(KEYINPUT86), .A3(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(G1971), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT86), .B1(new_n677), .B2(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n683));
  NAND2_X1  g258(.A1(G288), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT85), .A4(new_n570), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G16), .ZN(new_n687));
  OR2_X1    g262(.A1(G16), .A2(G23), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT33), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(G6), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G305), .B2(new_n676), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT32), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1981), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n682), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n681), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n677), .A2(KEYINPUT86), .A3(new_n678), .ZN(new_n698));
  OAI21_X1  g273(.A(G1971), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n675), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G24), .B(G290), .S(G16), .Z(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(G1986), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n490), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n492), .A2(G119), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n709));
  OAI221_X1 g284(.A(G2104), .B1(G107), .B2(new_n470), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n705), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n704), .B1(new_n712), .B2(new_n703), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n701), .A2(G1986), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n702), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n699), .A2(new_n682), .A3(new_n695), .A4(new_n691), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(KEYINPUT34), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n674), .B1(new_n700), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n696), .A2(new_n675), .A3(new_n699), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n722), .A2(new_n723), .A3(new_n718), .A4(new_n673), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n676), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n676), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n703), .A2(G32), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT95), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(G105), .B2(new_n474), .ZN(new_n736));
  AOI22_X1  g311(.A1(G129), .A2(new_n492), .B1(new_n490), .B2(G141), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n703), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n729), .B1(new_n739), .B2(new_n740), .C1(new_n746), .C2(G2084), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT98), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n495), .A2(G29), .A3(new_n496), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n703), .A2(G35), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT99), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n749), .B2(new_n751), .ZN(new_n754));
  OAI21_X1  g329(.A(G2090), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n746), .A2(G2084), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT93), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n727), .A2(new_n728), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n676), .A2(G21), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G286), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n620), .A2(new_n703), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(KEYINPUT96), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(KEYINPUT96), .B2(new_n765), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT88), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n597), .B2(new_n676), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1348), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n676), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT102), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n760), .A2(new_n767), .A3(new_n771), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  INV_X1    g353(.A(G127), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n481), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  NAND2_X1  g356(.A1(G103), .A2(G2104), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n780), .A2(G2105), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n490), .ZN(new_n786));
  INV_X1    g361(.A(G139), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G33), .B(new_n788), .S(G29), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2072), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n703), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n762), .B2(new_n763), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n703), .A2(G26), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT28), .Z(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT90), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n490), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n492), .A2(G128), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT91), .B(G2067), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n739), .B2(new_n740), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n703), .A2(G27), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G164), .B2(new_n703), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G19), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n813), .A2(KEYINPUT89), .A3(G16), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT89), .B1(new_n813), .B2(G16), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n814), .B(new_n815), .C1(new_n554), .C2(new_n676), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1341), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n806), .B2(new_n805), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n796), .A2(new_n808), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n753), .A2(new_n754), .A3(G2090), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n777), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AND4_X1   g396(.A1(new_n748), .A2(new_n756), .A3(new_n758), .A4(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n725), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n725), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(new_n725), .A2(new_n822), .ZN(G150));
  NAND2_X1  g402(.A1(new_n598), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n521), .ZN(new_n831));
  INV_X1    g406(.A(G55), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT104), .B(G93), .Z(new_n833));
  OAI22_X1  g408(.A1(new_n510), .A2(new_n832), .B1(new_n516), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n554), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n554), .A2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n829), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n835), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XOR2_X1   g422(.A(KEYINPUT107), .B(G37), .Z(new_n848));
  OAI211_X1 g423(.A(new_n785), .B(KEYINPUT106), .C1(new_n786), .C2(new_n787), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT105), .ZN(new_n850));
  INV_X1    g425(.A(G164), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n490), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n492), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n470), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n613), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n852), .A2(new_n853), .A3(new_n860), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n738), .B(new_n804), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n711), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n866), .ZN(new_n868));
  XNOR2_X1  g443(.A(G160), .B(new_n620), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G162), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n848), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g449(.A(G868), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n831), .B2(new_n834), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n598), .A2(G299), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n597), .A2(new_n602), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n879), .A2(KEYINPUT109), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(KEYINPUT108), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n597), .A2(new_n883), .A3(new_n602), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n884), .A3(new_n877), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n880), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT109), .B1(new_n879), .B2(new_n880), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n839), .B(new_n607), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n879), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n890), .B(KEYINPUT110), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(KEYINPUT110), .B2(new_n890), .ZN(new_n893));
  XNOR2_X1  g468(.A(G166), .B(G290), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n686), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT42), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n893), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n876), .B1(new_n898), .B2(new_n875), .ZN(G295));
  OAI21_X1  g474(.A(new_n876), .B1(new_n898), .B2(new_n875), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n901));
  AOI21_X1  g476(.A(G286), .B1(G171), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(G301), .A2(KEYINPUT111), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(G301), .A2(KEYINPUT111), .A3(G286), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n839), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n838), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT112), .A3(new_n909), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n906), .A2(KEYINPUT112), .A3(new_n838), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n891), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT113), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n891), .B2(KEYINPUT41), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n882), .A2(new_n877), .A3(KEYINPUT41), .A4(new_n884), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n879), .A2(KEYINPUT113), .A3(new_n880), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n908), .A2(new_n909), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n912), .B1(new_n919), .B2(KEYINPUT114), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT114), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n896), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n908), .A2(new_n879), .A3(new_n909), .ZN(new_n925));
  INV_X1    g500(.A(new_n888), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n910), .A2(new_n911), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n896), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n848), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  INV_X1    g506(.A(new_n896), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT43), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n929), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n924), .B1(new_n933), .B2(new_n928), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n503), .B2(new_n507), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n473), .A2(new_n475), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT71), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n473), .A2(KEYINPUT71), .A3(new_n475), .ZN(new_n948));
  INV_X1    g523(.A(G40), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n483), .B2(G2105), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n738), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n804), .B(G2067), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n714), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n712), .A2(new_n714), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n611), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n961));
  OAI21_X1  g536(.A(G40), .B1(new_n961), .B2(new_n470), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n476), .A2(new_n477), .A3(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT45), .B(new_n941), .C1(new_n503), .C2(new_n507), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n944), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n763), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(G2084), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n941), .C1(new_n503), .C2(new_n507), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n967), .A2(new_n963), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(G168), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n973));
  AND2_X1   g548(.A1(KEYINPUT121), .A2(G8), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n966), .A2(new_n971), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(G8), .A3(G286), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT122), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n972), .A2(new_n974), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT51), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT122), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n977), .A4(new_n975), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n577), .A2(new_n987), .A3(new_n578), .A4(new_n579), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n526), .A2(G61), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n521), .B1(new_n989), .B2(new_n575), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n578), .A2(new_n579), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n951), .B2(new_n942), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n684), .A2(G1976), .A3(new_n685), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(G8), .C1(new_n951), .C2(new_n942), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AND2_X1   g576(.A1(G288), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n997), .A2(new_n998), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT115), .B1(new_n1000), .B2(KEYINPUT52), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n965), .A2(new_n680), .ZN(new_n1012));
  INV_X1    g587(.A(G2090), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n967), .A2(new_n963), .A3(new_n1013), .A4(new_n970), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n528), .A2(new_n530), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1010), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1016), .B(KEYINPUT55), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n967), .A2(new_n963), .A3(new_n970), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1021), .A2(new_n1013), .B1(new_n965), .B2(new_n680), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT116), .B(new_n1020), .C1(new_n1022), .C2(new_n1011), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1009), .A2(new_n1019), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n944), .A2(new_n963), .A3(new_n811), .A4(new_n964), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n967), .A2(new_n963), .A3(new_n970), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n728), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1027), .A2(G2078), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n944), .A2(new_n963), .A3(new_n964), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1033), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT123), .B1(new_n1033), .B2(G171), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1025), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n986), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n986), .A2(new_n1037), .A3(KEYINPUT126), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n980), .A2(new_n985), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT62), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT127), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1046));
  AND4_X1   g621(.A1(new_n1040), .A2(new_n1041), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1011), .B(G286), .C1(new_n966), .C2(new_n971), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1000), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1049), .A2(new_n1024), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1052), .A2(new_n1053), .A3(new_n1048), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT63), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1056), .A2(new_n1057), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G288), .A2(G1976), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n997), .B2(new_n998), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n998), .B1(new_n1061), .B2(new_n988), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1024), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1009), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(G299), .B(KEYINPUT57), .Z(new_n1065));
  INV_X1    g640(.A(G1956), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1029), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n944), .A2(new_n963), .A3(new_n964), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1348), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n951), .A2(new_n942), .A3(G2067), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1072), .A2(new_n1029), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n963), .A2(new_n941), .A3(new_n851), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT118), .B1(new_n1076), .B2(G2067), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n598), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G299), .B(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1071), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n598), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(KEYINPUT60), .A3(new_n597), .A4(new_n1077), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1085), .A2(new_n1086), .B1(new_n1084), .B2(new_n1078), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT58), .B(G1341), .Z(new_n1089));
  OAI211_X1 g664(.A(new_n1088), .B(new_n1089), .C1(new_n951), .C2(new_n942), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n965), .B2(G1996), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1076), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n554), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT59), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n554), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1082), .A2(new_n1098), .A3(new_n1070), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1082), .B2(new_n1070), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1087), .B1(new_n1101), .B2(KEYINPUT120), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1097), .B(new_n1103), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1083), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n1033), .B2(G171), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n478), .A2(KEYINPUT124), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n961), .A2(KEYINPUT125), .ZN(new_n1108));
  OAI21_X1  g683(.A(G2105), .B1(new_n961), .B2(KEYINPUT125), .ZN(new_n1109));
  OAI211_X1 g684(.A(G40), .B(new_n1031), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n478), .A2(KEYINPUT124), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n944), .A3(new_n964), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1106), .B1(G171), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1025), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(G171), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1034), .A2(new_n1117), .A3(new_n1035), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n1042), .C1(KEYINPUT54), .C2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1059), .B(new_n1064), .C1(new_n1105), .C2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n960), .B1(new_n1047), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G290), .A2(G1986), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n952), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(KEYINPUT48), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1124), .A2(KEYINPUT48), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n958), .C2(new_n952), .ZN(new_n1127));
  INV_X1    g702(.A(new_n955), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n952), .B1(new_n1128), .B2(new_n738), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT46), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n952), .B2(new_n953), .ZN(new_n1131));
  NOR4_X1   g706(.A1(new_n944), .A2(new_n951), .A3(KEYINPUT46), .A4(G1996), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT47), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n954), .A2(new_n955), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1135), .A2(new_n956), .B1(G2067), .B2(new_n804), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1127), .B(new_n1134), .C1(new_n952), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1121), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g713(.A1(G401), .A2(new_n463), .A3(G227), .ZN(new_n1140));
  OAI21_X1  g714(.A(new_n1140), .B1(new_n670), .B2(new_n671), .ZN(new_n1141));
  INV_X1    g715(.A(new_n1141), .ZN(new_n1142));
  OAI211_X1 g716(.A(new_n873), .B(new_n1142), .C1(new_n937), .C2(new_n938), .ZN(G225));
  INV_X1    g717(.A(G225), .ZN(G308));
endmodule


