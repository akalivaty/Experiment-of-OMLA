//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(KEYINPUT65), .A3(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n199), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(G128), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n197), .A2(new_n198), .A3(new_n200), .A4(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n213), .A2(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n210), .A2(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n209), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n209), .A2(KEYINPUT81), .A3(new_n222), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT10), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT66), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT67), .A3(G131), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n236), .B2(new_n237), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n230), .A2(new_n232), .A3(new_n240), .A4(new_n233), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n201), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n246), .B(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n195), .B2(new_n200), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n245), .A2(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G101), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n256), .A3(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n195), .A2(new_n200), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n202), .A2(new_n203), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT68), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT68), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n208), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n222), .A3(KEYINPUT10), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n227), .A2(new_n244), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n244), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n224), .B(new_n221), .C1(new_n208), .C2(new_n205), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT81), .B1(new_n209), .B2(new_n222), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n258), .A2(new_n266), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n193), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n264), .A2(new_n208), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n225), .A2(new_n226), .B1(new_n278), .B2(new_n221), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n279), .B2(new_n269), .ZN(new_n280));
  OAI22_X1  g094(.A1(new_n271), .A2(new_n272), .B1(new_n265), .B2(new_n222), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT12), .A3(new_n244), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n274), .A3(new_n269), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT84), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n192), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n284), .B2(new_n192), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n276), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT83), .B(G469), .Z(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n275), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n284), .A3(new_n192), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n268), .B1(new_n282), .B2(new_n280), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n192), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT82), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT82), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n298), .B(new_n294), .C1(new_n295), .C2(new_n192), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n292), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n261), .A2(new_n262), .A3(new_n199), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n206), .A2(G143), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G122), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT91), .B1(new_n306), .B2(G116), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G122), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n305), .A2(new_n229), .B1(new_n313), .B2(new_n213), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n307), .A2(new_n310), .B1(G116), .B2(new_n306), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G107), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT92), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT13), .B1(new_n206), .B2(G143), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n199), .A3(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(KEYINPUT68), .A2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT68), .A2(G128), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(G143), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n317), .B1(new_n325), .B2(G134), .ZN(new_n326));
  AOI211_X1 g140(.A(KEYINPUT92), .B(new_n229), .C1(new_n321), .C2(new_n324), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n314), .B(new_n316), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n304), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(new_n229), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n229), .B1(new_n324), .B2(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT93), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n213), .B1(new_n312), .B2(KEYINPUT14), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n315), .B(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G134), .B1(new_n303), .B2(new_n304), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT93), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n330), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G217), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n187), .A2(new_n340), .A3(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT94), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n328), .A2(new_n339), .A3(KEYINPUT94), .A4(new_n341), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n328), .A2(new_n339), .ZN(new_n346));
  INV_X1    g160(.A(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT15), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G478), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n349), .A2(new_n290), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n349), .B2(new_n290), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT90), .B(G475), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(G125), .A3(G140), .ZN(new_n359));
  AOI21_X1  g173(.A(G140), .B1(new_n358), .B2(G125), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT75), .B(KEYINPUT16), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G125), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n362), .B1(new_n368), .B2(KEYINPUT74), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n358), .A2(G125), .A3(G140), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT75), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n194), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT16), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(G146), .A3(new_n361), .A4(new_n366), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n190), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n199), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n240), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT17), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(new_n199), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n240), .A3(new_n383), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n373), .A2(new_n378), .A3(new_n385), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT18), .A2(G131), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n381), .A2(new_n383), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT88), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n368), .A2(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n363), .A2(new_n397), .A3(new_n194), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n363), .A2(new_n397), .A3(KEYINPUT76), .A4(new_n194), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n369), .A2(G146), .A3(new_n370), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n402), .A2(new_n403), .B1(new_n384), .B2(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n392), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n210), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n392), .A2(new_n408), .A3(new_n405), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n357), .B1(new_n412), .B2(new_n290), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n392), .A2(new_n408), .A3(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n374), .A2(KEYINPUT19), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n363), .A2(new_n397), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n420), .A2(new_n194), .B1(new_n388), .B2(new_n390), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n396), .A2(new_n404), .B1(new_n421), .B2(new_n378), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n408), .B1(new_n422), .B2(KEYINPUT89), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n378), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n405), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n415), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n428), .A2(KEYINPUT20), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n405), .A2(new_n424), .A3(KEYINPUT89), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n409), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n422), .A2(KEYINPUT89), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n411), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n436), .B2(new_n429), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n414), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n355), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT85), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n190), .A2(G952), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G234), .B2(G237), .ZN(new_n443));
  INV_X1    g257(.A(G234), .ZN(new_n444));
  OAI211_X1 g258(.A(G902), .B(G953), .C1(new_n444), .C2(new_n379), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(G898), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT8), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT2), .B(G113), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G119), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT5), .ZN(new_n455));
  INV_X1    g269(.A(G119), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(G116), .ZN(new_n457));
  INV_X1    g271(.A(new_n453), .ZN(new_n458));
  OAI211_X1 g272(.A(G113), .B(new_n457), .C1(new_n458), .C2(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n222), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n222), .B1(new_n454), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n450), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n451), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n454), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n255), .A2(new_n465), .A3(new_n257), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n460), .A3(new_n449), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n278), .A2(new_n368), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n249), .A2(new_n251), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n201), .B2(new_n246), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G125), .ZN(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(new_n472), .B2(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n463), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n471), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n468), .A2(new_n471), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n472), .A2(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n466), .A2(new_n460), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  INV_X1    g301(.A(new_n449), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT6), .A3(new_n467), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n481), .A2(new_n492), .A3(new_n494), .ZN(new_n497));
  AOI211_X1 g311(.A(new_n441), .B(new_n448), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  AND4_X1   g312(.A1(new_n188), .A2(new_n302), .A3(new_n439), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n382), .A2(G210), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT27), .Z(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT26), .B(G101), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n243), .B1(new_n238), .B2(G131), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n506), .B(new_n240), .C1(new_n236), .C2(new_n237), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n252), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n229), .A2(G137), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n231), .A2(G134), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n242), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n265), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n465), .B(KEYINPUT70), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n465), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n508), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT28), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n513), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n244), .B2(new_n252), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n514), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n504), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT69), .B(KEYINPUT30), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n508), .A2(new_n513), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n508), .B2(new_n513), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n465), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n504), .A3(new_n521), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n508), .A2(new_n513), .A3(new_n525), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n520), .B2(new_n529), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n515), .B1(new_n536), .B2(new_n465), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n504), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT71), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n524), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT31), .B1(new_n537), .B2(new_n504), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT11), .B1(new_n231), .B2(G134), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT66), .B1(new_n546), .B2(new_n232), .ZN(new_n547));
  INV_X1    g361(.A(new_n237), .ZN(new_n548));
  OAI21_X1  g362(.A(G131), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n243), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n470), .B1(new_n551), .B2(new_n239), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n528), .B1(new_n552), .B2(new_n519), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n516), .B1(new_n553), .B2(new_n535), .ZN(new_n554));
  NOR4_X1   g368(.A1(new_n554), .A2(new_n533), .A3(new_n503), .A4(new_n515), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n543), .B1(new_n544), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT71), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n540), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT32), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n542), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n523), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n522), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n520), .B(new_n514), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n504), .A2(KEYINPUT29), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n290), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n531), .A2(new_n521), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n503), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n518), .A2(new_n504), .A3(new_n523), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G472), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n560), .A2(new_n561), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G217), .B1(new_n444), .B2(G902), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT73), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n373), .A2(new_n378), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n261), .A2(new_n262), .A3(new_n456), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n206), .A2(G119), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT24), .B(G110), .ZN(new_n584));
  OR3_X1    g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT23), .B1(new_n206), .B2(G119), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n456), .B2(G128), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n322), .A2(KEYINPUT23), .A3(G119), .A4(new_n323), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n581), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n594));
  INV_X1    g408(.A(G110), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n594), .A2(new_n596), .B1(new_n400), .B2(new_n401), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n378), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n591), .B1(new_n373), .B2(new_n378), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n378), .A2(new_n597), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT25), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n607), .B2(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n608), .B(KEYINPUT25), .C1(new_n607), .C2(KEYINPUT77), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n580), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n603), .A2(new_n606), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT79), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n579), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT80), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n613), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n499), .A2(new_n577), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  INV_X1    g443(.A(new_n188), .ZN(new_n630));
  INV_X1    g444(.A(new_n299), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n279), .A2(new_n277), .A3(new_n269), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT12), .B1(new_n281), .B2(new_n244), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n284), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n193), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n298), .B1(new_n635), .B2(new_n294), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n290), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G469), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n630), .B1(new_n638), .B2(new_n292), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n539), .B2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n542), .A2(new_n640), .A3(new_n558), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(new_n627), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n498), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT20), .B1(new_n428), .B2(new_n430), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n436), .A2(new_n432), .A3(new_n429), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n413), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n348), .A2(KEYINPUT33), .A3(new_n342), .ZN(new_n648));
  INV_X1    g462(.A(G478), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(G902), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n349), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n349), .B2(new_n652), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n648), .B(new_n650), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n349), .A2(new_n290), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n649), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n647), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n644), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n643), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NOR2_X1   g478(.A1(new_n438), .A2(new_n354), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n498), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n643), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n593), .A2(new_n598), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n621), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n613), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n499), .A2(new_n642), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT98), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NOR2_X1   g495(.A1(KEYINPUT99), .A2(G900), .ZN(new_n682));
  AND2_X1   g496(.A1(KEYINPUT99), .A2(G900), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n446), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n443), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n681), .B1(new_n665), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n441), .B1(new_n496), .B2(new_n497), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n613), .B2(new_n674), .ZN(new_n689));
  INV_X1    g503(.A(new_n686), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n438), .A2(new_n354), .A3(KEYINPUT100), .A4(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n577), .A2(new_n692), .A3(new_n639), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n577), .A2(new_n692), .A3(new_n639), .A4(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  INV_X1    g512(.A(new_n532), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n503), .B2(new_n566), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n560), .A2(new_n561), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT102), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n686), .B(KEYINPUT39), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n639), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n496), .A2(new_n497), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT38), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n355), .A2(new_n438), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n711), .A2(new_n676), .A3(new_n441), .A4(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n705), .A2(new_n708), .A3(new_n709), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n658), .A2(new_n716), .A3(new_n688), .A4(new_n686), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n655), .A2(new_n657), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n688), .A3(new_n438), .A4(new_n686), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n675), .B1(new_n719), .B2(KEYINPUT103), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n577), .A2(new_n639), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n676), .A3(new_n717), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n577), .A4(new_n639), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  NAND2_X1  g542(.A1(new_n289), .A2(new_n290), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT105), .A3(G469), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n284), .A2(new_n192), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT84), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n283), .A3(new_n286), .ZN(new_n734));
  AOI21_X1  g548(.A(G902), .B1(new_n734), .B2(new_n276), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(new_n735), .B2(new_n301), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n188), .A2(new_n730), .A3(new_n736), .A4(new_n292), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n661), .A2(new_n577), .A3(new_n627), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT106), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT41), .B(G113), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n577), .A2(new_n627), .A3(new_n666), .A4(new_n737), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NAND3_X1  g557(.A1(new_n676), .A2(new_n439), .A3(new_n498), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n730), .A2(new_n736), .A3(new_n188), .A4(new_n292), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n577), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  INV_X1    g562(.A(new_n448), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n688), .A2(new_n438), .A3(new_n355), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n563), .A2(new_n564), .B1(new_n566), .B2(KEYINPUT28), .ZN(new_n752));
  OAI22_X1  g566(.A1(new_n544), .A2(new_n555), .B1(new_n752), .B2(new_n504), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n540), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n640), .A2(new_n754), .A3(new_n623), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n758), .A2(new_n718), .A3(new_n438), .A4(new_n686), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n658), .B2(new_n686), .ZN(new_n760));
  INV_X1    g574(.A(new_n688), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n745), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n640), .A2(new_n754), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT107), .B1(new_n763), .B2(new_n675), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n676), .A2(new_n754), .A3(new_n765), .A4(new_n640), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  NOR2_X1   g583(.A1(new_n759), .A2(new_n760), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n710), .A2(new_n441), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n188), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n732), .A2(new_n275), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n634), .B2(new_n193), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n774), .B2(G902), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n292), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT109), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n292), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n772), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n577), .A2(new_n770), .A3(new_n780), .A4(new_n627), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n559), .B1(new_n539), .B2(new_n541), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n576), .A2(new_n561), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(new_n623), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n770), .A4(new_n780), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT110), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  NAND2_X1  g607(.A1(new_n665), .A2(new_n686), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n795));
  INV_X1    g609(.A(new_n691), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT111), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n687), .B2(new_n691), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n577), .A3(new_n627), .A4(new_n780), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  AOI21_X1  g616(.A(new_n438), .B1(new_n657), .B2(new_n655), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT43), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n438), .B2(KEYINPUT113), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT114), .B1(new_n806), .B2(new_n807), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n641), .B(new_n676), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT44), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n771), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(KEYINPUT115), .B(new_n771), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n301), .A2(new_n290), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n297), .B2(new_n299), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  OAI21_X1  g635(.A(G469), .B1(new_n296), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT46), .B(new_n819), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT112), .A3(new_n292), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n820), .A2(new_n822), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n818), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(KEYINPUT46), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT112), .B1(new_n823), .B2(new_n292), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n188), .B(new_n706), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n813), .B2(new_n812), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(new_n817), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  OAI21_X1  g646(.A(new_n188), .B1(new_n827), .B2(new_n828), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT47), .B(new_n188), .C1(new_n827), .C2(new_n828), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n627), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n658), .A3(new_n686), .A4(new_n771), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n577), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NAND2_X1  g656(.A1(new_n808), .A2(new_n443), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n730), .A2(new_n736), .A3(new_n292), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(new_n772), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n786), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT48), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n838), .A2(new_n845), .A3(new_n685), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n659), .A2(new_n660), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n704), .A4(new_n703), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n685), .B1(new_n806), .B2(new_n807), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n755), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n761), .A3(new_n745), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n442), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n848), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT118), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n848), .A2(new_n858), .A3(new_n851), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n711), .A2(new_n441), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n852), .A3(new_n737), .A4(new_n755), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT50), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n718), .A2(new_n438), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n704), .A2(new_n849), .A3(new_n703), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n846), .A2(new_n767), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n771), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n853), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n844), .A2(new_n188), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n837), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n867), .B2(new_n871), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n860), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n860), .B(new_n877), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n767), .A2(new_n770), .A3(new_n780), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n771), .A2(new_n439), .A3(new_n686), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n771), .A2(new_n439), .A3(KEYINPUT117), .A4(new_n686), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n675), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n577), .A3(new_n639), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n801), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n789), .A2(new_n791), .A3(new_n887), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n746), .A2(new_n577), .B1(new_n751), .B2(new_n755), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(new_n738), .A3(new_n742), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n889), .A2(new_n892), .A3(new_n738), .A4(new_n742), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n658), .A2(new_n665), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n644), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n639), .A2(new_n627), .A3(new_n642), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n628), .A2(new_n677), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n676), .A2(new_n630), .A3(new_n690), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n761), .A2(new_n712), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n777), .A2(new_n779), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n702), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n727), .A2(new_n697), .A3(new_n768), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n695), .A2(new_n696), .B1(new_n767), .B2(new_n762), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT52), .A3(new_n727), .A4(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  AND4_X1   g724(.A1(KEYINPUT53), .A2(new_n628), .A3(new_n677), .A4(new_n896), .ZN(new_n911));
  INV_X1    g725(.A(new_n890), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n887), .A3(new_n912), .A4(new_n788), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n906), .B2(new_n908), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(KEYINPUT54), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n899), .A2(new_n909), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT54), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n879), .A2(new_n921), .B1(G952), .B2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n844), .B(KEYINPUT49), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n630), .A2(new_n441), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n711), .A2(new_n623), .A3(new_n803), .A4(new_n924), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n705), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(G75));
  OAI211_X1 g741(.A(G210), .B(G902), .C1(new_n910), .C2(new_n914), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n491), .A2(new_n489), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n484), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT122), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n190), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n928), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n928), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n929), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n942), .B2(new_n933), .ZN(G51));
  XOR2_X1   g757(.A(new_n818), .B(KEYINPUT123), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT57), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT54), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n917), .A2(new_n918), .ZN(new_n947));
  INV_X1    g761(.A(new_n914), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n945), .B1(new_n949), .B2(new_n915), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n289), .ZN(new_n951));
  OAI211_X1 g765(.A(G902), .B(new_n825), .C1(new_n910), .C2(new_n914), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n936), .B1(new_n951), .B2(new_n953), .ZN(G54));
  AND2_X1   g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  OAI211_X1 g769(.A(G902), .B(new_n955), .C1(new_n910), .C2(new_n914), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n956), .A2(KEYINPUT125), .A3(new_n428), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT125), .B1(new_n956), .B2(new_n428), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n936), .B1(new_n956), .B2(new_n428), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  OAI21_X1  g774(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n921), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n962), .B(new_n965), .C1(new_n949), .C2(new_n915), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n937), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n910), .B2(new_n914), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n619), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n673), .B(KEYINPUT126), .Z(new_n974));
  OAI211_X1 g788(.A(new_n971), .B(new_n974), .C1(new_n910), .C2(new_n914), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n937), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n937), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  NAND2_X1  g794(.A1(G224), .A2(G953), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n898), .A2(G953), .B1(new_n447), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n930), .B1(G898), .B2(new_n190), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  AOI21_X1  g798(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n536), .B(new_n420), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n907), .A2(new_n727), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n714), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n707), .A2(new_n868), .A3(new_n894), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n577), .A3(new_n627), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n831), .A2(new_n841), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n988), .B1(new_n997), .B2(new_n190), .ZN(new_n998));
  INV_X1    g812(.A(new_n988), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n829), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n901), .A3(new_n786), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n792), .A2(new_n801), .A3(new_n989), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n831), .A2(new_n841), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1001), .B1(new_n1006), .B2(new_n190), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n986), .B(new_n987), .C1(new_n998), .C2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n990), .B(KEYINPUT62), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(new_n995), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n999), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1007), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT127), .A4(new_n985), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1008), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  INV_X1    g830(.A(new_n1006), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n898), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n571), .A2(new_n504), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n936), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1016), .B1(new_n997), .B2(new_n898), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1021), .A2(new_n504), .A3(new_n571), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n572), .A2(new_n532), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1016), .B(new_n1023), .C1(new_n919), .C2(new_n910), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(G57));
endmodule


