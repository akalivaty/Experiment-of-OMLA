

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595;

  XNOR2_X1 U328 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U329 ( .A(n397), .B(n396), .ZN(n565) );
  XOR2_X1 U330 ( .A(n344), .B(n343), .Z(n533) );
  XNOR2_X1 U331 ( .A(n432), .B(KEYINPUT48), .ZN(n433) );
  INV_X1 U332 ( .A(KEYINPUT95), .ZN(n336) );
  XNOR2_X1 U333 ( .A(n384), .B(KEYINPUT9), .ZN(n385) );
  XNOR2_X1 U334 ( .A(n434), .B(n433), .ZN(n544) );
  XNOR2_X1 U335 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n486) );
  XNOR2_X1 U336 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U337 ( .A(n386), .B(n385), .ZN(n389) );
  XNOR2_X1 U338 ( .A(n487), .B(n486), .ZN(n527) );
  XNOR2_X1 U339 ( .A(n395), .B(n394), .ZN(n396) );
  INV_X1 U340 ( .A(G183GAT), .ZN(n465) );
  NOR2_X1 U341 ( .A1(n543), .A2(n463), .ZN(n575) );
  XNOR2_X1 U342 ( .A(n381), .B(n380), .ZN(n583) );
  INV_X1 U343 ( .A(KEYINPUT104), .ZN(n491) );
  XNOR2_X1 U344 ( .A(n465), .B(KEYINPUT124), .ZN(n466) );
  XNOR2_X1 U345 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U346 ( .A(n467), .B(n466), .ZN(G1350GAT) );
  XNOR2_X1 U347 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(G15GAT), .B(G127GAT), .Z(n404) );
  XOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT0), .Z(n441) );
  XNOR2_X1 U350 ( .A(n404), .B(n441), .ZN(n297) );
  XNOR2_X1 U351 ( .A(G71GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n296), .B(G120GAT), .ZN(n355) );
  XNOR2_X1 U353 ( .A(n297), .B(n355), .ZN(n302) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n298), .B(G134GAT), .ZN(n391) );
  XOR2_X1 U356 ( .A(KEYINPUT20), .B(n391), .Z(n300) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U359 ( .A(n302), .B(n301), .Z(n311) );
  XNOR2_X1 U360 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n303), .B(KEYINPUT17), .ZN(n304) );
  XOR2_X1 U362 ( .A(n304), .B(KEYINPUT19), .Z(n306) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n342) );
  XOR2_X1 U365 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n308) );
  XNOR2_X1 U366 ( .A(G99GAT), .B(KEYINPUT84), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n342), .B(n309), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n543) );
  XOR2_X1 U370 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n313) );
  XOR2_X1 U371 ( .A(G50GAT), .B(G162GAT), .Z(n387) );
  XOR2_X1 U372 ( .A(G22GAT), .B(G155GAT), .Z(n403) );
  XNOR2_X1 U373 ( .A(n387), .B(n403), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U375 ( .A(n314), .B(G106GAT), .Z(n320) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n315), .B(KEYINPUT2), .ZN(n445) );
  XOR2_X1 U378 ( .A(n445), .B(G211GAT), .Z(n317) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n318), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U383 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n322) );
  XNOR2_X1 U384 ( .A(KEYINPUT88), .B(KEYINPUT90), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U386 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G148GAT), .Z(n326) );
  XNOR2_X1 U388 ( .A(KEYINPUT70), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U389 ( .A(n326), .B(n325), .ZN(n347) );
  XNOR2_X1 U390 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n327), .B(KEYINPUT21), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n347), .B(n335), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n479) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G204GAT), .Z(n331) );
  XNOR2_X1 U395 ( .A(G190GAT), .B(G176GAT), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n341) );
  XNOR2_X1 U397 ( .A(G8GAT), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n332), .B(KEYINPUT77), .ZN(n398) );
  XOR2_X1 U399 ( .A(G36GAT), .B(G218GAT), .Z(n383) );
  XOR2_X1 U400 ( .A(n398), .B(n383), .Z(n334) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U402 ( .A(n334), .B(n333), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n335), .B(G64GAT), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n344) );
  INV_X1 U405 ( .A(n342), .ZN(n343) );
  INV_X1 U406 ( .A(n533), .ZN(n435) );
  XOR2_X1 U407 ( .A(G85GAT), .B(G92GAT), .Z(n346) );
  XNOR2_X1 U408 ( .A(G99GAT), .B(G106GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n390) );
  XNOR2_X1 U410 ( .A(n347), .B(n390), .ZN(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n349) );
  XNOR2_X1 U412 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n351) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n357) );
  XNOR2_X1 U418 ( .A(G64GAT), .B(G57GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n354), .B(KEYINPUT13), .ZN(n402) );
  XNOR2_X1 U420 ( .A(n355), .B(n402), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n586) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G197GAT), .Z(n361) );
  XNOR2_X1 U424 ( .A(G169GAT), .B(G141GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U426 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n363) );
  XNOR2_X1 U427 ( .A(G113GAT), .B(G8GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT67), .B(G1GAT), .Z(n412) );
  XOR2_X1 U431 ( .A(G22GAT), .B(G50GAT), .Z(n367) );
  XNOR2_X1 U432 ( .A(G43GAT), .B(G36GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U434 ( .A(n412), .B(n368), .Z(n370) );
  NAND2_X1 U435 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U437 ( .A(n371), .B(KEYINPUT65), .Z(n379) );
  INV_X1 U438 ( .A(KEYINPUT8), .ZN(n372) );
  NAND2_X1 U439 ( .A1(G29GAT), .A2(n372), .ZN(n375) );
  INV_X1 U440 ( .A(G29GAT), .ZN(n373) );
  NAND2_X1 U441 ( .A1(n373), .A2(KEYINPUT8), .ZN(n374) );
  NAND2_X1 U442 ( .A1(n375), .A2(n374), .ZN(n377) );
  XNOR2_X1 U443 ( .A(KEYINPUT7), .B(KEYINPUT66), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n382), .B(KEYINPUT29), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n386) );
  AND2_X1 U448 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X1 U449 ( .A(n387), .B(KEYINPUT73), .Z(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U452 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n393) );
  XNOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT75), .ZN(n392) );
  XOR2_X1 U454 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U455 ( .A(KEYINPUT76), .B(n565), .ZN(n574) );
  XNOR2_X1 U456 ( .A(n574), .B(KEYINPUT36), .ZN(n484) );
  XOR2_X1 U457 ( .A(KEYINPUT14), .B(n398), .Z(n400) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U460 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n418) );
  XOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n410) );
  XNOR2_X1 U467 ( .A(G71GAT), .B(KEYINPUT15), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n411), .B(G78GAT), .Z(n414) );
  XNOR2_X1 U470 ( .A(n412), .B(G183GAT), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U472 ( .A(n416), .B(n415), .Z(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n591) );
  NAND2_X1 U474 ( .A1(n484), .A2(n591), .ZN(n420) );
  XOR2_X1 U475 ( .A(KEYINPUT45), .B(KEYINPUT117), .Z(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  NOR2_X1 U477 ( .A1(n583), .A2(n421), .ZN(n422) );
  NAND2_X1 U478 ( .A1(n586), .A2(n422), .ZN(n431) );
  XNOR2_X1 U479 ( .A(n586), .B(KEYINPUT41), .ZN(n569) );
  NAND2_X1 U480 ( .A1(n583), .A2(n569), .ZN(n425) );
  XOR2_X1 U481 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT114), .B(n423), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(KEYINPUT113), .B(n591), .ZN(n551) );
  NAND2_X1 U485 ( .A1(n426), .A2(n551), .ZN(n427) );
  NOR2_X1 U486 ( .A1(n565), .A2(n427), .ZN(n429) );
  XNOR2_X1 U487 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n430) );
  NAND2_X1 U489 ( .A1(n431), .A2(n430), .ZN(n434) );
  XNOR2_X1 U490 ( .A(KEYINPUT64), .B(KEYINPUT118), .ZN(n432) );
  NAND2_X1 U491 ( .A1(n435), .A2(n544), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n436), .B(KEYINPUT121), .ZN(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT54), .B(n437), .ZN(n460) );
  XOR2_X1 U494 ( .A(G85GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U497 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U500 ( .A(n444), .B(KEYINPUT4), .Z(n447) );
  XNOR2_X1 U501 ( .A(n445), .B(KEYINPUT5), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U503 ( .A(KEYINPUT74), .B(G155GAT), .Z(n449) );
  XNOR2_X1 U504 ( .A(G127GAT), .B(G148GAT), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U506 ( .A(n451), .B(n450), .Z(n459) );
  XOR2_X1 U507 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT6), .B(KEYINPUT92), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT94), .B(G57GAT), .Z(n455) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(G120GAT), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n530) );
  NAND2_X1 U515 ( .A1(n460), .A2(n530), .ZN(n582) );
  NOR2_X1 U516 ( .A1(n479), .A2(n582), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U519 ( .A(n575), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n464), .A2(n551), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n543), .A2(n533), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n479), .A2(n468), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT25), .ZN(n474) );
  XOR2_X1 U524 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n471) );
  NAND2_X1 U525 ( .A1(n479), .A2(n543), .ZN(n470) );
  XOR2_X1 U526 ( .A(n471), .B(n470), .Z(n581) );
  XNOR2_X1 U527 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(n533), .ZN(n477) );
  OR2_X1 U529 ( .A1(n581), .A2(n477), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n530), .A2(n475), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT99), .ZN(n482) );
  NOR2_X1 U533 ( .A1(n530), .A2(n477), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT97), .B(n478), .Z(n558) );
  XOR2_X1 U535 ( .A(n479), .B(KEYINPUT28), .Z(n539) );
  NAND2_X1 U536 ( .A1(n558), .A2(n539), .ZN(n542) );
  XNOR2_X1 U537 ( .A(n543), .B(KEYINPUT87), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n542), .A2(n480), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n499), .A2(n591), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT102), .B(n483), .ZN(n485) );
  NAND2_X1 U542 ( .A1(n485), .A2(n484), .ZN(n487) );
  NAND2_X1 U543 ( .A1(n583), .A2(n586), .ZN(n495) );
  NOR2_X1 U544 ( .A1(n527), .A2(n495), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n488), .Z(n513) );
  NOR2_X1 U546 ( .A1(n543), .A2(n513), .ZN(n494) );
  XOR2_X1 U547 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n490) );
  XNOR2_X1 U548 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n492) );
  INV_X1 U550 ( .A(n495), .ZN(n500) );
  INV_X1 U551 ( .A(n591), .ZN(n496) );
  NOR2_X1 U552 ( .A1(n496), .A2(n574), .ZN(n497) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n497), .Z(n498) );
  NOR2_X1 U554 ( .A1(n499), .A2(n498), .ZN(n516) );
  NAND2_X1 U555 ( .A1(n500), .A2(n516), .ZN(n507) );
  NOR2_X1 U556 ( .A1(n530), .A2(n507), .ZN(n501) );
  XOR2_X1 U557 ( .A(G1GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U558 ( .A(KEYINPUT34), .B(n502), .ZN(G1324GAT) );
  NOR2_X1 U559 ( .A1(n533), .A2(n507), .ZN(n503) );
  XOR2_X1 U560 ( .A(G8GAT), .B(n503), .Z(G1325GAT) );
  NOR2_X1 U561 ( .A1(n543), .A2(n507), .ZN(n505) );
  XNOR2_X1 U562 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  NOR2_X1 U565 ( .A1(n539), .A2(n507), .ZN(n508) );
  XOR2_X1 U566 ( .A(G22GAT), .B(n508), .Z(G1327GAT) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n509), .B(KEYINPUT39), .ZN(n511) );
  NOR2_X1 U569 ( .A1(n530), .A2(n513), .ZN(n510) );
  XOR2_X1 U570 ( .A(n511), .B(n510), .Z(G1328GAT) );
  NOR2_X1 U571 ( .A1(n533), .A2(n513), .ZN(n512) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U573 ( .A1(n539), .A2(n513), .ZN(n514) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  INV_X1 U575 ( .A(n583), .ZN(n515) );
  NAND2_X1 U576 ( .A1(n515), .A2(n569), .ZN(n528) );
  INV_X1 U577 ( .A(n528), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n517), .A2(n516), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n530), .A2(n522), .ZN(n518) );
  XOR2_X1 U580 ( .A(n518), .B(KEYINPUT42), .Z(n519) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NOR2_X1 U582 ( .A1(n533), .A2(n522), .ZN(n520) );
  XOR2_X1 U583 ( .A(G64GAT), .B(n520), .Z(G1333GAT) );
  NOR2_X1 U584 ( .A1(n543), .A2(n522), .ZN(n521) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n539), .ZN(n526) );
  XOR2_X1 U587 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n524) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(KEYINPUT109), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n530), .A2(n538), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT110), .B(n531), .Z(n532) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n538), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n543), .A2(n538), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT112), .B(n536), .Z(n537) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(n537), .ZN(G1338GAT) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U603 ( .A(KEYINPUT44), .B(n540), .Z(n541) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT119), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n554), .A2(n583), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U611 ( .A1(n554), .A2(n569), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  INV_X1 U613 ( .A(n554), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n552), .Z(n553) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U618 ( .A1(n554), .A2(n574), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U621 ( .A1(n544), .A2(n558), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n581), .A2(n559), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n583), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U626 ( .A1(n566), .A2(n569), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U629 ( .A1(n591), .A2(n566), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n575), .A2(n583), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n571) );
  NAND2_X1 U636 ( .A1(n575), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT123), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT60), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(n580), .Z(n585) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n593) );
  NAND2_X1 U648 ( .A1(n593), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n589) );
  INV_X1 U651 ( .A(n586), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n593), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G204GAT), .B(n590), .Z(G1353GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n593), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U657 ( .A1(n593), .A2(n484), .ZN(n594) );
  XNOR2_X1 U658 ( .A(n594), .B(KEYINPUT62), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

