

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576;

  XOR2_X1 U319 ( .A(G1GAT), .B(G127GAT), .Z(n354) );
  XNOR2_X1 U320 ( .A(n371), .B(n370), .ZN(n372) );
  INV_X1 U321 ( .A(G92GAT), .ZN(n377) );
  XOR2_X1 U322 ( .A(n309), .B(n308), .Z(n553) );
  XNOR2_X1 U323 ( .A(KEYINPUT101), .B(n468), .ZN(n515) );
  XOR2_X1 U324 ( .A(KEYINPUT77), .B(KEYINPUT13), .Z(n287) );
  AND2_X1 U325 ( .A1(G230GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U326 ( .A(KEYINPUT114), .B(KEYINPUT45), .ZN(n365) );
  XNOR2_X1 U327 ( .A(n366), .B(n365), .ZN(n383) );
  NOR2_X1 U328 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U329 ( .A(n369), .B(n288), .ZN(n370) );
  XNOR2_X1 U330 ( .A(n334), .B(n436), .ZN(n338) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G57GAT), .Z(n376) );
  XNOR2_X1 U332 ( .A(n338), .B(n337), .ZN(n339) );
  INV_X1 U333 ( .A(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U334 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U335 ( .A1(n487), .A2(n489), .ZN(n491) );
  XNOR2_X1 U336 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U337 ( .A(KEYINPUT84), .B(n553), .ZN(n540) );
  XNOR2_X1 U338 ( .A(n568), .B(n406), .ZN(n556) );
  XOR2_X1 U339 ( .A(KEYINPUT38), .B(n493), .Z(n501) );
  XOR2_X1 U340 ( .A(n463), .B(KEYINPUT28), .Z(n528) );
  XNOR2_X1 U341 ( .A(n449), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U342 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n290) );
  XNOR2_X1 U344 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n289) );
  XNOR2_X1 U345 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U346 ( .A(n291), .B(KEYINPUT82), .Z(n293) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G106GAT), .Z(n369) );
  XNOR2_X1 U348 ( .A(n369), .B(KEYINPUT9), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U350 ( .A(G92GAT), .B(KEYINPUT83), .Z(n295) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n417) );
  XNOR2_X1 U353 ( .A(n417), .B(KEYINPUT81), .ZN(n297) );
  AND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U357 ( .A(G162GAT), .B(KEYINPUT80), .Z(n301) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(G218GAT), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n323) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n302), .B(G85GAT), .ZN(n340) );
  XNOR2_X1 U362 ( .A(n323), .B(n340), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U364 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U365 ( .A(KEYINPUT73), .B(G43GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U367 ( .A(KEYINPUT72), .B(n307), .ZN(n388) );
  INV_X1 U368 ( .A(n388), .ZN(n308) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(KEYINPUT95), .Z(n311) );
  XNOR2_X1 U370 ( .A(KEYINPUT2), .B(KEYINPUT94), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n312), .B(G155GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n344) );
  XOR2_X1 U375 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n316) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n344), .B(n317), .ZN(n327) );
  XOR2_X1 U379 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n319) );
  NAND2_X1 U380 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n322) );
  XOR2_X1 U382 ( .A(G204GAT), .B(G211GAT), .Z(n321) );
  XNOR2_X1 U383 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n420) );
  XOR2_X1 U385 ( .A(n322), .B(n420), .Z(n325) );
  XNOR2_X1 U386 ( .A(G22GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n463) );
  XOR2_X1 U389 ( .A(KEYINPUT1), .B(KEYINPUT96), .Z(n329) );
  XNOR2_X1 U390 ( .A(G162GAT), .B(KEYINPUT6), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U392 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n331) );
  XNOR2_X1 U393 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U396 ( .A(G113GAT), .B(KEYINPUT0), .Z(n436) );
  XOR2_X1 U397 ( .A(n354), .B(n376), .Z(n336) );
  NAND2_X1 U398 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U400 ( .A(n339), .B(KEYINPUT99), .Z(n342) );
  XNOR2_X1 U401 ( .A(n340), .B(KEYINPUT98), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n468) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT87), .Z(n346) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n351) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n287), .B(n347), .ZN(n371) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G183GAT), .Z(n414) );
  XOR2_X1 U410 ( .A(n371), .B(n414), .Z(n349) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n364) );
  XOR2_X1 U414 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n353) );
  XNOR2_X1 U415 ( .A(G57GAT), .B(G64GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n355) );
  XOR2_X1 U417 ( .A(n355), .B(n354), .Z(n357) );
  XNOR2_X1 U418 ( .A(G155GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U420 ( .A(n358), .B(KEYINPUT88), .Z(n362) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n360) );
  XNOR2_X1 U422 ( .A(G22GAT), .B(G15GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n387) );
  XNOR2_X1 U424 ( .A(n387), .B(KEYINPUT89), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U426 ( .A(n364), .B(n363), .Z(n473) );
  INV_X1 U427 ( .A(n473), .ZN(n571) );
  XNOR2_X1 U428 ( .A(KEYINPUT36), .B(n540), .ZN(n487) );
  NOR2_X1 U429 ( .A1(n571), .A2(n487), .ZN(n366) );
  XOR2_X1 U430 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n368) );
  XNOR2_X1 U431 ( .A(G148GAT), .B(G204GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U433 ( .A(n372), .B(KEYINPUT33), .Z(n375) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G64GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT78), .ZN(n419) );
  XNOR2_X1 U436 ( .A(n419), .B(KEYINPUT79), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n380) );
  XNOR2_X1 U438 ( .A(G85GAT), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n568) );
  NAND2_X1 U440 ( .A1(n383), .A2(n568), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT115), .ZN(n405) );
  XOR2_X1 U442 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n386) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(G8GAT), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n390) );
  XOR2_X1 U446 ( .A(n388), .B(n387), .Z(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n404) );
  NAND2_X1 U449 ( .A1(G229GAT), .A2(G233GAT), .ZN(n398) );
  XOR2_X1 U450 ( .A(G113GAT), .B(G141GAT), .Z(n394) );
  XNOR2_X1 U451 ( .A(G50GAT), .B(G197GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U453 ( .A(G36GAT), .B(G29GAT), .Z(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT76), .B(G1GAT), .Z(n400) );
  XNOR2_X1 U457 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U460 ( .A(n404), .B(n403), .Z(n503) );
  INV_X1 U461 ( .A(n503), .ZN(n564) );
  NAND2_X1 U462 ( .A1(n405), .A2(n564), .ZN(n412) );
  NAND2_X1 U463 ( .A1(n553), .A2(n571), .ZN(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n406) );
  NOR2_X1 U465 ( .A1(n564), .A2(n556), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n407), .B(KEYINPUT46), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n410), .B(KEYINPUT47), .ZN(n411) );
  NAND2_X1 U468 ( .A1(n412), .A2(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(KEYINPUT48), .B(n413), .Z(n526) );
  XOR2_X1 U470 ( .A(G218GAT), .B(n414), .Z(n416) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U473 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U476 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n424) );
  XNOR2_X1 U477 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(G169GAT), .B(n425), .Z(n443) );
  XOR2_X1 U480 ( .A(n426), .B(n443), .Z(n456) );
  NOR2_X1 U481 ( .A1(n526), .A2(n456), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  NOR2_X1 U483 ( .A1(n515), .A2(n429), .ZN(n563) );
  NAND2_X1 U484 ( .A1(n463), .A2(n563), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n430), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U486 ( .A(G127GAT), .B(G120GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G15GAT), .B(G183GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n447) );
  XOR2_X1 U489 ( .A(G176GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U490 ( .A(G99GAT), .B(G190GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U492 ( .A(n435), .B(G134GAT), .Z(n438) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT66), .Z(n440) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U498 ( .A(n442), .B(n441), .Z(n445) );
  XNOR2_X1 U499 ( .A(n443), .B(KEYINPUT91), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(n447), .B(n446), .Z(n459) );
  INV_X1 U502 ( .A(n459), .ZN(n530) );
  NAND2_X1 U503 ( .A1(n448), .A2(n530), .ZN(n452) );
  NOR2_X1 U504 ( .A1(n540), .A2(n452), .ZN(n451) );
  XNOR2_X1 U505 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n449) );
  NOR2_X1 U506 ( .A1(n571), .A2(n452), .ZN(n455) );
  INV_X1 U507 ( .A(G183GAT), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(KEYINPUT124), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n479) );
  INV_X1 U511 ( .A(n456), .ZN(n518) );
  XNOR2_X1 U512 ( .A(n518), .B(KEYINPUT102), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n457), .ZN(n465) );
  NAND2_X1 U514 ( .A1(n465), .A2(n515), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT103), .B(n458), .Z(n525) );
  NOR2_X1 U516 ( .A1(n528), .A2(n525), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n460), .A2(n459), .ZN(n471) );
  NAND2_X1 U518 ( .A1(n530), .A2(n518), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n463), .A2(n461), .ZN(n462) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n462), .Z(n467) );
  NOR2_X1 U521 ( .A1(n530), .A2(n463), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT26), .ZN(n562) );
  NAND2_X1 U523 ( .A1(n562), .A2(n465), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT104), .B(n472), .ZN(n488) );
  XOR2_X1 U528 ( .A(KEYINPUT90), .B(KEYINPUT16), .Z(n475) );
  NAND2_X1 U529 ( .A1(n473), .A2(n540), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  AND2_X1 U531 ( .A1(n488), .A2(n476), .ZN(n504) );
  AND2_X1 U532 ( .A1(n503), .A2(n568), .ZN(n492) );
  NAND2_X1 U533 ( .A1(n504), .A2(n492), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT105), .ZN(n485) );
  NAND2_X1 U535 ( .A1(n515), .A2(n485), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n518), .A2(n485), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT106), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT35), .B(KEYINPUT107), .Z(n483) );
  NAND2_X1 U541 ( .A1(n485), .A2(n530), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n484), .Z(G1326GAT) );
  NAND2_X1 U544 ( .A1(n485), .A2(n528), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U547 ( .A1(n571), .A2(n488), .ZN(n489) );
  XOR2_X1 U548 ( .A(KEYINPUT108), .B(KEYINPUT37), .Z(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n513) );
  NAND2_X1 U550 ( .A1(n513), .A2(n492), .ZN(n493) );
  NAND2_X1 U551 ( .A1(n515), .A2(n501), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n496), .Z(G1328GAT) );
  NAND2_X1 U554 ( .A1(n501), .A2(n518), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT110), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n501), .A2(n530), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT40), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n501), .A2(n528), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U562 ( .A1(n556), .A2(n503), .ZN(n514) );
  AND2_X1 U563 ( .A1(n504), .A2(n514), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n515), .A2(n510), .ZN(n505) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n505), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U567 ( .A(G64GAT), .B(KEYINPUT111), .Z(n508) );
  NAND2_X1 U568 ( .A1(n510), .A2(n518), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n508), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n530), .A2(n510), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U573 ( .A1(n510), .A2(n528), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  AND2_X1 U575 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U579 ( .A1(n518), .A2(n522), .ZN(n519) );
  XNOR2_X1 U580 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U581 ( .A(G99GAT), .B(KEYINPUT113), .Z(n521) );
  NAND2_X1 U582 ( .A1(n522), .A2(n530), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n528), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U588 ( .A(KEYINPUT116), .B(n527), .ZN(n544) );
  INV_X1 U589 ( .A(n544), .ZN(n529) );
  NOR2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n539) );
  NOR2_X1 U592 ( .A1(n564), .A2(n539), .ZN(n533) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  NOR2_X1 U595 ( .A1(n556), .A2(n539), .ZN(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n571), .A2(n539), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NAND2_X1 U606 ( .A1(n562), .A2(n544), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n564), .A2(n552), .ZN(n545) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n556), .A2(n552), .ZN(n550) );
  XOR2_X1 U610 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT120), .B(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n571), .A2(n552), .ZN(n551) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n564), .A2(n452), .ZN(n555) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n555), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n452), .A2(n556), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n574) );
  NOR2_X1 U628 ( .A1(n564), .A2(n574), .ZN(n566) );
  XNOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n568), .A2(n574), .ZN(n570) );
  XNOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n574), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(n572), .Z(n573) );
  XNOR2_X1 U637 ( .A(G211GAT), .B(n573), .ZN(G1354GAT) );
  NOR2_X1 U638 ( .A1(n487), .A2(n574), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT62), .B(n575), .Z(n576) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(n576), .ZN(G1355GAT) );
endmodule

