//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT80), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n205), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(KEYINPUT14), .ZN(new_n209));
  NOR3_X1   g008(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n209), .A2(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT15), .B1(new_n213), .B2(G43gat), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G50gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n206), .A2(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n214), .B2(new_n216), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(G50gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT81), .A4(KEYINPUT15), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT82), .B1(new_n215), .B2(G50gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(new_n216), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n215), .A2(KEYINPUT82), .A3(G50gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT15), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n212), .A2(new_n218), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G15gat), .B(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(G1gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT16), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n235), .B(new_n236), .C1(G1gat), .C2(new_n232), .ZN(new_n237));
  INV_X1    g036(.A(G15gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G22gat), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G15gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n234), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(G1gat), .B1(new_n239), .B2(new_n241), .ZN(new_n243));
  OAI21_X1  g042(.A(G8gat), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n202), .B1(new_n231), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n237), .A2(new_n244), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n219), .B1(new_n210), .B2(KEYINPUT80), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n206), .A2(new_n207), .ZN(new_n249));
  OAI22_X1  g048(.A1(new_n248), .A2(new_n249), .B1(new_n204), .B2(new_n205), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n217), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n223), .A3(new_n229), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(new_n225), .A3(new_n222), .A4(new_n220), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n247), .A2(KEYINPUT83), .A3(new_n251), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n231), .A2(new_n245), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n246), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G229gat), .A2(G233gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT13), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT84), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT17), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n231), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n251), .A3(KEYINPUT17), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n247), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n261), .A3(new_n259), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT18), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n260), .A2(new_n272), .A3(new_n262), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n268), .A2(KEYINPUT18), .A3(new_n261), .A4(new_n259), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n264), .A2(new_n271), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G113gat), .B(G141gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G197gat), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT11), .B(G169gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT12), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n273), .A3(new_n274), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT85), .A3(new_n270), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n280), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT85), .B1(new_n269), .B2(new_n270), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(KEYINPUT23), .B2(new_n292), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n294), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT24), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n304), .B2(new_n303), .ZN(new_n306));
  AND3_X1   g105(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n290), .B1(new_n302), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n309), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n315));
  OR2_X1    g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  OR3_X1    g116(.A1(new_n298), .A2(new_n292), .A3(KEYINPUT26), .ZN(new_n318));
  INV_X1    g117(.A(new_n303), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(KEYINPUT26), .B2(new_n292), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n310), .B1(KEYINPUT24), .B2(new_n319), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(new_n290), .A3(new_n299), .A4(new_n301), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n312), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT1), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  OAI221_X1 g129(.A(new_n328), .B1(new_n326), .B2(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n331), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n312), .A2(new_n324), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n331), .B(new_n332), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n335), .A2(G227gat), .A3(G233gat), .A4(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G15gat), .B(G43gat), .Z(new_n342));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n335), .A2(new_n338), .ZN(new_n347));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT34), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT34), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n345), .A2(new_n350), .A3(new_n352), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n354), .B2(new_n357), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(KEYINPUT22), .B2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G211gat), .B(G218gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G141gat), .B(G148gat), .Z(new_n369));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(KEYINPUT72), .B(G155gat), .Z(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT73), .B(G162gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n372), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n368), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(new_n368), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT29), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT31), .B(G50gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n240), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n240), .B2(new_n391), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n388), .B(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n361), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(KEYINPUT35), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT70), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G226gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n336), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n325), .A2(new_n381), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n407), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n368), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT69), .B1(new_n409), .B2(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n407), .ZN(new_n413));
  INV_X1    g212(.A(new_n408), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n415), .B2(KEYINPUT69), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n403), .B(new_n411), .C1(new_n416), .C2(new_n368), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT71), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n411), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n410), .B2(new_n421), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n423), .B2(new_n384), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT30), .A4(new_n403), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n384), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n403), .B1(new_n428), .B2(new_n411), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n418), .B2(new_n417), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  INV_X1    g232(.A(new_n379), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n334), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n380), .A2(new_n438), .A3(new_n337), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n434), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT74), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n337), .A2(new_n379), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n435), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n447), .B2(new_n443), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n448), .ZN(new_n450));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT0), .ZN(new_n452));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n449), .B2(new_n450), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n433), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n449), .A2(new_n450), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n454), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT77), .A3(new_n457), .A4(new_n456), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n398), .A2(new_n432), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n458), .B2(new_n459), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n464), .A2(KEYINPUT75), .A3(new_n457), .A4(new_n456), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n462), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n427), .A3(new_n430), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT35), .B1(new_n472), .B2(new_n397), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n441), .A2(new_n443), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(KEYINPUT39), .C1(new_n443), .C2(new_n447), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n454), .C1(KEYINPUT39), .C2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT40), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n479), .A2(new_n480), .A3(new_n461), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n431), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n428), .A2(new_n483), .A3(new_n411), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n402), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n424), .A2(new_n483), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT38), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n423), .B2(new_n384), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n368), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n410), .A2(KEYINPUT79), .A3(new_n368), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT79), .B1(new_n410), .B2(new_n368), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(KEYINPUT37), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n484), .A2(new_n495), .A3(new_n402), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n487), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n460), .A2(new_n465), .A3(new_n462), .A4(new_n417), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n482), .B(new_n396), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n359), .B2(new_n360), .ZN(new_n501));
  INV_X1    g300(.A(new_n360), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT36), .A3(new_n358), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n472), .A2(new_n395), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n289), .B1(new_n474), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G190gat), .B(G218gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(KEYINPUT90), .A2(G99gat), .A3(G106gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(KEYINPUT8), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT7), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G85gat), .ZN(new_n518));
  INV_X1    g317(.A(G92gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n513), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n512), .A2(new_n517), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G99gat), .B(G106gat), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n508), .B2(new_n509), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n527), .A2(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n528));
  INV_X1    g327(.A(new_n524), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n522), .A4(new_n517), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n266), .A2(new_n267), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n231), .A2(new_n265), .B1(new_n530), .B2(new_n525), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT91), .A3(new_n267), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n525), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n231), .ZN(new_n539));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT92), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n546), .B(new_n543), .C1(new_n534), .C2(new_n536), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n507), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  AND4_X1   g347(.A1(KEYINPUT91), .A2(new_n266), .A3(new_n267), .A4(new_n531), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT91), .B1(new_n535), .B2(new_n267), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n546), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n553));
  INV_X1    g352(.A(new_n507), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT87), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G134gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G162gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n548), .A2(new_n555), .A3(KEYINPUT88), .A4(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(G57gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT9), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT86), .B1(new_n565), .B2(G57gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(G64gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n576), .A3(new_n566), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n571), .B1(new_n570), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n569), .A2(new_n572), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G127gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n247), .B1(new_n582), .B2(new_n581), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G155gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n564), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n525), .A2(new_n580), .A3(new_n530), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n531), .A2(new_n581), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT93), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n600), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n531), .A2(KEYINPUT93), .A3(new_n581), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n602), .B1(new_n607), .B2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(G230gat), .A2(G233gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n599), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n600), .A2(new_n604), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n580), .B1(new_n525), .B2(new_n530), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n606), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n601), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n619));
  INV_X1    g418(.A(new_n602), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT10), .B1(new_n605), .B2(new_n606), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT94), .B1(new_n622), .B2(new_n602), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n623), .A3(new_n609), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n612), .A2(new_n599), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n613), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n595), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n506), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n471), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n233), .ZN(G1324gat));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n631), .A2(KEYINPUT96), .A3(new_n432), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT96), .B1(new_n631), .B2(new_n432), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(G8gat), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n631), .A2(new_n432), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT16), .B(G8gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n635), .B2(new_n636), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(KEYINPUT42), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n634), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n637), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n646), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(G1325gat));
  INV_X1    g451(.A(new_n631), .ZN(new_n653));
  AOI21_X1  g452(.A(G15gat), .B1(new_n653), .B2(new_n361), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT100), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n501), .A2(new_n503), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n631), .A2(new_n238), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n395), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n594), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n562), .A2(new_n563), .ZN(new_n664));
  INV_X1    g463(.A(new_n613), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n624), .A2(new_n626), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT95), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND4_X1   g468(.A1(new_n506), .A2(new_n663), .A3(new_n664), .A4(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n471), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n204), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n674), .B(new_n564), .C1(new_n474), .C2(new_n505), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n499), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT103), .B1(new_n499), .B2(new_n504), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n474), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n664), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n679), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n669), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT102), .B1(new_n283), .B2(new_n288), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n286), .A2(new_n287), .ZN(new_n683));
  INV_X1    g482(.A(new_n284), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(new_n282), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n680), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n678), .B2(new_n664), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  INV_X1    g491(.A(new_n689), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n691), .A2(new_n692), .A3(new_n675), .A4(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n690), .A2(new_n694), .A3(new_n471), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n673), .B1(new_n695), .B2(new_n204), .ZN(G1328gat));
  AOI21_X1  g495(.A(G36gat), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n670), .A2(new_n431), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n690), .A2(new_n694), .A3(new_n432), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n205), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT106), .B(new_n700), .C1(new_n701), .C2(new_n205), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n670), .A2(new_n215), .A3(new_n361), .ZN(new_n707));
  INV_X1    g506(.A(new_n680), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n656), .A3(new_n693), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT47), .B(new_n707), .C1(new_n709), .C2(new_n215), .ZN(new_n710));
  INV_X1    g509(.A(new_n707), .ZN(new_n711));
  INV_X1    g510(.A(new_n690), .ZN(new_n712));
  INV_X1    g511(.A(new_n656), .ZN(new_n713));
  INV_X1    g512(.A(new_n694), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n715), .B2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n716), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g516(.A1(new_n396), .A2(G50gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n670), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n708), .A2(new_n396), .A3(new_n693), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT48), .B(new_n719), .C1(new_n720), .C2(new_n213), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n712), .A2(new_n395), .A3(new_n714), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(G50gat), .B1(new_n670), .B2(new_n718), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g523(.A(new_n688), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n595), .A2(new_n725), .A3(new_n669), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n678), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n671), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n730), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n432), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n727), .B(KEYINPUT107), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n737), .A3(new_n733), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n736), .A2(G71gat), .A3(new_n713), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n727), .A2(new_n361), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(G71gat), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n395), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT109), .B(G78gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  INV_X1    g547(.A(new_n679), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n725), .A2(new_n594), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n629), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n671), .A2(new_n518), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n750), .A2(new_n629), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n708), .A2(new_n471), .A3(new_n758), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n756), .A2(new_n757), .B1(new_n518), .B2(new_n759), .ZN(G1336gat));
  INV_X1    g559(.A(new_n754), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n749), .B2(new_n750), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n431), .A2(new_n519), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n763), .A2(new_n669), .A3(new_n764), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n708), .A2(new_n432), .A3(new_n758), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n519), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT52), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  OAI221_X1 g568(.A(new_n769), .B1(new_n766), .B2(new_n519), .C1(new_n756), .C2(new_n764), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(G1337gat));
  INV_X1    g570(.A(new_n758), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n680), .A2(new_n713), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n680), .A2(KEYINPUT110), .A3(new_n713), .A4(new_n772), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(G99gat), .A3(new_n776), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n359), .A2(new_n360), .A3(G99gat), .A4(new_n669), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT111), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n763), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n777), .B(KEYINPUT112), .C1(new_n763), .C2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n396), .A2(G106gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n629), .B(new_n786), .C1(new_n761), .C2(new_n762), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n680), .A2(new_n395), .A3(new_n772), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(KEYINPUT53), .A3(G106gat), .ZN(new_n789));
  OR2_X1    g588(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n793), .A2(new_n794), .B1(new_n787), .B2(KEYINPUT113), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n260), .A2(new_n262), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n261), .B1(new_n268), .B2(new_n259), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n279), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(KEYINPUT115), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n288), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n629), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n667), .A2(new_n668), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n618), .A2(new_n620), .A3(new_n610), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n618), .A2(new_n620), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n610), .B1(new_n809), .B2(KEYINPUT94), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n621), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n609), .C1(new_n622), .C2(new_n602), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n599), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n806), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n608), .B2(new_n610), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n624), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n805), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n804), .B1(new_n819), .B2(new_n688), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n564), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n667), .A2(new_n668), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n664), .A2(new_n803), .A3(new_n822), .A4(new_n815), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n594), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n595), .A2(new_n725), .A3(new_n629), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT116), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n802), .A2(new_n801), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n685), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n819), .A2(new_n564), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n564), .B2(new_n820), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n827), .B(new_n828), .C1(new_n832), .C2(new_n594), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(new_n396), .A3(new_n361), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n431), .A2(new_n471), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n326), .A3(new_n289), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n725), .A3(new_n836), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n326), .B2(new_n839), .ZN(G1340gat));
  NOR2_X1   g639(.A1(new_n837), .A2(new_n669), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(new_n327), .ZN(G1341gat));
  NOR2_X1   g641(.A1(new_n837), .A2(new_n663), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(new_n586), .ZN(G1342gat));
  NOR2_X1   g643(.A1(new_n431), .A2(new_n564), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n471), .A2(G134gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n835), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT56), .Z(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n837), .B2(new_n564), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n395), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(new_n289), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n624), .A2(new_n816), .ZN(new_n854));
  INV_X1    g653(.A(new_n814), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT119), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n817), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n822), .B(new_n853), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n669), .B2(new_n830), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n629), .A2(KEYINPUT117), .A3(new_n803), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n564), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n594), .B1(new_n867), .B2(new_n823), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(new_n825), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n396), .A2(new_n852), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n851), .A2(new_n852), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n836), .A2(new_n656), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n289), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n851), .A2(new_n872), .ZN(new_n877));
  INV_X1    g676(.A(G141gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n878), .A3(new_n853), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n879), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n873), .A2(new_n725), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(new_n876), .ZN(G1344gat));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n629), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n826), .A2(new_n833), .A3(new_n870), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n664), .A2(new_n890), .A3(new_n822), .A4(new_n815), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT121), .B1(new_n819), .B2(new_n564), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n803), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n594), .B1(new_n867), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n595), .A2(new_n853), .A3(new_n629), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n395), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n888), .A2(new_n889), .B1(new_n896), .B2(new_n852), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n826), .A2(new_n833), .A3(KEYINPUT120), .A4(new_n870), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n669), .B(new_n872), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n885), .B1(new_n899), .B2(KEYINPUT122), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n887), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g701(.A(KEYINPUT59), .B(new_n885), .C1(new_n873), .C2(new_n629), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n886), .B1(new_n902), .B2(new_n903), .ZN(G1345gat));
  OAI21_X1  g703(.A(new_n375), .B1(new_n874), .B2(new_n663), .ZN(new_n905));
  INV_X1    g704(.A(new_n375), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n877), .A2(new_n906), .A3(new_n594), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1346gat));
  OAI21_X1  g707(.A(new_n376), .B1(new_n874), .B2(new_n564), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n713), .A2(new_n376), .A3(new_n471), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n845), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n851), .B2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n432), .A2(new_n671), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n835), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(G169gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(new_n289), .ZN(new_n916));
  INV_X1    g715(.A(new_n914), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n725), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(G1348gat));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n629), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g720(.A(new_n308), .B1(new_n914), .B2(new_n663), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(new_n594), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n313), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n914), .B2(new_n564), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n926), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(KEYINPUT61), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n926), .B2(KEYINPUT61), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n927), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n309), .A3(new_n664), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1351gat));
  NOR4_X1   g734(.A1(new_n713), .A2(new_n671), .A3(new_n432), .A4(new_n396), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n834), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n725), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n913), .A2(new_n656), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n897), .B2(new_n898), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n853), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  NOR3_X1   g742(.A1(new_n937), .A2(G204gat), .A3(new_n669), .ZN(new_n944));
  XNOR2_X1  g743(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n941), .ZN(new_n947));
  OAI21_X1  g746(.A(G204gat), .B1(new_n947), .B2(new_n669), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1353gat));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n888), .A2(new_n889), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n896), .A2(new_n852), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n898), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954));
  INV_X1    g753(.A(new_n940), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n953), .A2(new_n954), .A3(new_n594), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n941), .B2(new_n594), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n953), .A2(new_n594), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n956), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n938), .A2(new_n363), .A3(new_n594), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1354gat));
  OAI21_X1  g768(.A(G218gat), .B1(new_n947), .B2(new_n564), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n938), .A2(new_n364), .A3(new_n664), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1355gat));
endmodule


