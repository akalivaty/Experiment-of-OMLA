

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U556 ( .A1(n606), .A2(n524), .ZN(n621) );
  INV_X1 U557 ( .A(G651), .ZN(n530) );
  INV_X1 U558 ( .A(G2104), .ZN(n546) );
  AND2_X1 U559 ( .A1(n602), .A2(n601), .ZN(G164) );
  XNOR2_X1 U560 ( .A(n549), .B(n548), .ZN(n892) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n732) );
  BUF_X1 U562 ( .A(n607), .Z(n532) );
  BUF_X1 U563 ( .A(n892), .Z(n522) );
  AND2_X1 U564 ( .A1(n547), .A2(n546), .ZN(n549) );
  NOR2_X1 U565 ( .A1(n621), .A2(n976), .ZN(n623) );
  AND2_X1 U566 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U567 ( .A1(n732), .A2(n603), .ZN(n631) );
  AND2_X1 U568 ( .A1(n991), .A2(n528), .ZN(n703) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n548) );
  NOR2_X2 U570 ( .A1(n547), .A2(n546), .ZN(n888) );
  INV_X1 U571 ( .A(KEYINPUT73), .ZN(n619) );
  NOR2_X1 U572 ( .A1(n631), .A2(n604), .ZN(n605) );
  OR2_X1 U573 ( .A1(n638), .A2(n986), .ZN(n635) );
  AND2_X1 U574 ( .A1(n525), .A2(n755), .ZN(n523) );
  AND2_X1 U575 ( .A1(n631), .A2(G1341), .ZN(n524) );
  AND2_X1 U576 ( .A1(n736), .A2(n735), .ZN(n525) );
  INV_X2 U577 ( .A(G2105), .ZN(n547) );
  OR2_X1 U578 ( .A1(n713), .A2(n712), .ZN(n526) );
  AND2_X1 U579 ( .A1(n710), .A2(n709), .ZN(n527) );
  OR2_X1 U580 ( .A1(n713), .A2(n702), .ZN(n528) );
  INV_X1 U581 ( .A(KEYINPUT64), .ZN(n622) );
  INV_X1 U582 ( .A(KEYINPUT101), .ZN(n636) );
  INV_X1 U583 ( .A(n631), .ZN(n660) );
  INV_X1 U584 ( .A(KEYINPUT29), .ZN(n658) );
  INV_X1 U585 ( .A(KEYINPUT103), .ZN(n687) );
  XNOR2_X1 U586 ( .A(n683), .B(KEYINPUT32), .ZN(n693) );
  BUF_X1 U587 ( .A(n631), .Z(n676) );
  INV_X1 U588 ( .A(G543), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n531), .B(KEYINPUT65), .ZN(n607) );
  NAND2_X1 U591 ( .A1(G160), .A2(G40), .ZN(n731) );
  AND2_X1 U592 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U593 ( .A1(G2105), .A2(n546), .ZN(n596) );
  NOR2_X1 U594 ( .A1(G651), .A2(n577), .ZN(n797) );
  XOR2_X1 U595 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NOR2_X1 U596 ( .A1(n556), .A2(n555), .ZN(G160) );
  XNOR2_X1 U597 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n532), .A2(G89), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT4), .ZN(n535) );
  NOR2_X4 U600 ( .A1(n577), .A2(n530), .ZN(n792) );
  NAND2_X1 U601 ( .A1(G76), .A2(n792), .ZN(n534) );
  NAND2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT5), .ZN(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n541) );
  NOR2_X1 U605 ( .A1(G543), .A2(n530), .ZN(n537) );
  XOR2_X1 U606 ( .A(KEYINPUT1), .B(n537), .Z(n612) );
  BUF_X1 U607 ( .A(n612), .Z(n796) );
  NAND2_X1 U608 ( .A1(G63), .A2(n796), .ZN(n539) );
  NAND2_X1 U609 ( .A1(G51), .A2(n797), .ZN(n538) );
  NAND2_X1 U610 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G168) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U615 ( .A1(n892), .A2(G137), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G101), .A2(n596), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT23), .B(n550), .Z(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G113), .A2(n888), .ZN(n554) );
  NOR2_X2 U620 ( .A1(G2104), .A2(n547), .ZN(n889) );
  NAND2_X1 U621 ( .A1(G125), .A2(n889), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G64), .A2(n796), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G52), .A2(n797), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT66), .B(n559), .Z(n566) );
  NAND2_X1 U627 ( .A1(n532), .A2(G90), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT67), .B(n560), .Z(n562) );
  NAND2_X1 U629 ( .A1(n792), .A2(G77), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U631 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(n567), .ZN(G171) );
  NAND2_X1 U635 ( .A1(G88), .A2(n532), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G75), .A2(n792), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G62), .A2(n796), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G50), .A2(n797), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(G166) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  NAND2_X1 U643 ( .A1(G49), .A2(n797), .ZN(n575) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n796), .A2(n576), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n577), .A2(G87), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U649 ( .A1(G86), .A2(n532), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G61), .A2(n796), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G73), .A2(n792), .ZN(n582) );
  XNOR2_X1 U653 ( .A(n582), .B(KEYINPUT85), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n583), .B(KEYINPUT2), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n797), .A2(G48), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U658 ( .A1(G85), .A2(n532), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G72), .A2(n792), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U661 ( .A1(G60), .A2(n796), .ZN(n591) );
  NAND2_X1 U662 ( .A1(G47), .A2(n797), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  OR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(G290) );
  AND2_X1 U665 ( .A1(G138), .A2(n892), .ZN(n595) );
  INV_X1 U666 ( .A(KEYINPUT90), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n595), .B(n594), .ZN(n602) );
  AND2_X1 U668 ( .A1(n889), .A2(G126), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G114), .A2(n888), .ZN(n598) );
  BUF_X2 U670 ( .A(n596), .Z(n894) );
  NAND2_X1 U671 ( .A1(G102), .A2(n894), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  INV_X1 U674 ( .A(n731), .ZN(n603) );
  INV_X1 U675 ( .A(G1996), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT26), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(G81), .ZN(n608) );
  XNOR2_X1 U678 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G68), .A2(n792), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n611), .B(KEYINPUT13), .ZN(n615) );
  NAND2_X1 U682 ( .A1(n612), .A2(G56), .ZN(n613) );
  XNOR2_X1 U683 ( .A(KEYINPUT14), .B(n613), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n616), .B(KEYINPUT72), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G43), .A2(n797), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n618), .A2(n617), .ZN(n620) );
  XNOR2_X2 U687 ( .A(n620), .B(n619), .ZN(n976) );
  XNOR2_X1 U688 ( .A(n623), .B(n622), .ZN(n638) );
  NAND2_X1 U689 ( .A1(G92), .A2(n532), .ZN(n625) );
  NAND2_X1 U690 ( .A1(G79), .A2(n792), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U692 ( .A1(G66), .A2(n796), .ZN(n627) );
  NAND2_X1 U693 ( .A1(G54), .A2(n797), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U696 ( .A(KEYINPUT15), .B(n630), .Z(n916) );
  INV_X1 U697 ( .A(n916), .ZN(n986) );
  NOR2_X1 U698 ( .A1(n660), .A2(G1348), .ZN(n633) );
  NOR2_X1 U699 ( .A1(G2067), .A2(n676), .ZN(n632) );
  NOR2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n637), .B(n636), .ZN(n640) );
  NAND2_X1 U703 ( .A1(n638), .A2(n986), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U705 ( .A(n641), .B(KEYINPUT102), .ZN(n653) );
  NAND2_X1 U706 ( .A1(n660), .A2(G2072), .ZN(n642) );
  XNOR2_X1 U707 ( .A(KEYINPUT27), .B(n642), .ZN(n645) );
  NAND2_X1 U708 ( .A1(G1956), .A2(n676), .ZN(n643) );
  XOR2_X1 U709 ( .A(KEYINPUT100), .B(n643), .Z(n644) );
  NOR2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n654) );
  NAND2_X1 U711 ( .A1(G65), .A2(n796), .ZN(n647) );
  NAND2_X1 U712 ( .A1(G53), .A2(n797), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U714 ( .A1(G91), .A2(n532), .ZN(n649) );
  NAND2_X1 U715 ( .A1(G78), .A2(n792), .ZN(n648) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n981) );
  NAND2_X1 U718 ( .A1(n654), .A2(n981), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U720 ( .A1(n654), .A2(n981), .ZN(n655) );
  XOR2_X1 U721 ( .A(n655), .B(KEYINPUT28), .Z(n656) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n659), .B(n658), .ZN(n666) );
  NOR2_X1 U724 ( .A1(n660), .A2(G1961), .ZN(n661) );
  XOR2_X1 U725 ( .A(KEYINPUT98), .B(n661), .Z(n664) );
  XOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .Z(n957) );
  NOR2_X1 U727 ( .A1(n957), .A2(n676), .ZN(n662) );
  XNOR2_X1 U728 ( .A(KEYINPUT99), .B(n662), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n670) );
  NAND2_X1 U730 ( .A1(n670), .A2(G171), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n675) );
  NOR2_X1 U732 ( .A1(G2084), .A2(n676), .ZN(n689) );
  NAND2_X1 U733 ( .A1(G8), .A2(n676), .ZN(n713) );
  NOR2_X1 U734 ( .A1(G1966), .A2(n713), .ZN(n684) );
  NOR2_X1 U735 ( .A1(n689), .A2(n684), .ZN(n667) );
  NAND2_X1 U736 ( .A1(G8), .A2(n667), .ZN(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT30), .B(n668), .ZN(n669) );
  NOR2_X1 U738 ( .A1(G168), .A2(n669), .ZN(n672) );
  NOR2_X1 U739 ( .A1(G171), .A2(n670), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U741 ( .A(KEYINPUT31), .B(n673), .Z(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n686), .A2(G286), .ZN(n681) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n713), .ZN(n678) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n676), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n679), .A2(G303), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n682), .A2(G8), .ZN(n683) );
  INV_X1 U750 ( .A(n684), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n688), .B(n687), .ZN(n691) );
  NAND2_X1 U752 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U755 ( .A(n694), .B(KEYINPUT104), .ZN(n706) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n701) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n701), .A2(n695), .ZN(n982) );
  AND2_X1 U759 ( .A1(n706), .A2(n982), .ZN(n698) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U761 ( .A(n713), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n980), .A2(n696), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U764 ( .A1(n699), .A2(KEYINPUT33), .ZN(n700) );
  INV_X1 U765 ( .A(n700), .ZN(n704) );
  XOR2_X1 U766 ( .A(G1981), .B(G305), .Z(n991) );
  NAND2_X1 U767 ( .A1(n701), .A2(KEYINPUT33), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n710) );
  NOR2_X1 U769 ( .A1(G2090), .A2(G303), .ZN(n705) );
  NAND2_X1 U770 ( .A1(G8), .A2(n705), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n708), .A2(n713), .ZN(n709) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n711) );
  XOR2_X1 U774 ( .A(n711), .B(KEYINPUT24), .Z(n712) );
  NAND2_X1 U775 ( .A1(n527), .A2(n526), .ZN(n748) );
  NAND2_X1 U776 ( .A1(G119), .A2(n889), .ZN(n715) );
  NAND2_X1 U777 ( .A1(G131), .A2(n522), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U779 ( .A1(G107), .A2(n888), .ZN(n717) );
  NAND2_X1 U780 ( .A1(G95), .A2(n894), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n907) );
  NAND2_X1 U783 ( .A1(G1991), .A2(n907), .ZN(n729) );
  NAND2_X1 U784 ( .A1(G117), .A2(n888), .ZN(n721) );
  NAND2_X1 U785 ( .A1(G129), .A2(n889), .ZN(n720) );
  NAND2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n894), .A2(G105), .ZN(n722) );
  XOR2_X1 U788 ( .A(KEYINPUT38), .B(n722), .Z(n723) );
  NOR2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U790 ( .A(n725), .B(KEYINPUT94), .ZN(n727) );
  NAND2_X1 U791 ( .A1(G141), .A2(n522), .ZN(n726) );
  NAND2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n911) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n911), .ZN(n728) );
  NAND2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U795 ( .A(KEYINPUT95), .B(n730), .ZN(n948) );
  NOR2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n760) );
  XOR2_X1 U797 ( .A(n760), .B(KEYINPUT96), .Z(n733) );
  NOR2_X1 U798 ( .A1(n948), .A2(n733), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n752), .B(KEYINPUT97), .ZN(n736) );
  XNOR2_X1 U800 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U801 ( .A1(n988), .A2(n760), .ZN(n734) );
  XOR2_X1 U802 ( .A(KEYINPUT91), .B(n734), .Z(n735) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n757) );
  NAND2_X1 U804 ( .A1(G116), .A2(n888), .ZN(n738) );
  NAND2_X1 U805 ( .A1(G128), .A2(n889), .ZN(n737) );
  NAND2_X1 U806 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U807 ( .A(KEYINPUT35), .B(n739), .Z(n746) );
  XNOR2_X1 U808 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n740) );
  XNOR2_X1 U809 ( .A(n740), .B(KEYINPUT34), .ZN(n744) );
  NAND2_X1 U810 ( .A1(G104), .A2(n894), .ZN(n742) );
  NAND2_X1 U811 ( .A1(G140), .A2(n522), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U813 ( .A(n744), .B(n743), .Z(n745) );
  NOR2_X1 U814 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n747), .ZN(n900) );
  NOR2_X1 U816 ( .A1(n757), .A2(n900), .ZN(n939) );
  NAND2_X1 U817 ( .A1(n760), .A2(n939), .ZN(n755) );
  NAND2_X1 U818 ( .A1(n748), .A2(n523), .ZN(n762) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n911), .ZN(n943) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n907), .ZN(n938) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n749) );
  NOR2_X1 U822 ( .A1(n938), .A2(n749), .ZN(n750) );
  XOR2_X1 U823 ( .A(KEYINPUT105), .B(n750), .Z(n751) );
  NOR2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U825 ( .A1(n943), .A2(n753), .ZN(n754) );
  XNOR2_X1 U826 ( .A(KEYINPUT39), .B(n754), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n757), .A2(n900), .ZN(n933) );
  NAND2_X1 U829 ( .A1(n758), .A2(n933), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U832 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G860), .ZN(n803) );
  OR2_X1 U835 ( .A1(n976), .A2(n803), .ZN(G153) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U839 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U840 ( .A(G223), .B(KEYINPUT71), .ZN(n833) );
  NAND2_X1 U841 ( .A1(n833), .A2(G567), .ZN(n766) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  NAND2_X1 U844 ( .A1(G301), .A2(G868), .ZN(n767) );
  XNOR2_X1 U845 ( .A(n767), .B(KEYINPUT74), .ZN(n769) );
  INV_X1 U846 ( .A(G868), .ZN(n815) );
  NAND2_X1 U847 ( .A1(n815), .A2(n986), .ZN(n768) );
  NAND2_X1 U848 ( .A1(n769), .A2(n768), .ZN(G284) );
  NOR2_X1 U849 ( .A1(G286), .A2(n815), .ZN(n770) );
  XNOR2_X1 U850 ( .A(n770), .B(KEYINPUT77), .ZN(n772) );
  NAND2_X1 U851 ( .A1(n981), .A2(n815), .ZN(n771) );
  NAND2_X1 U852 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U853 ( .A(KEYINPUT78), .B(n773), .Z(G297) );
  NAND2_X1 U854 ( .A1(n803), .A2(G559), .ZN(n774) );
  NAND2_X1 U855 ( .A1(n774), .A2(n916), .ZN(n775) );
  XNOR2_X1 U856 ( .A(n775), .B(KEYINPUT80), .ZN(n777) );
  XOR2_X1 U857 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n776) );
  XNOR2_X1 U858 ( .A(n777), .B(n776), .ZN(G148) );
  OR2_X1 U859 ( .A1(G559), .A2(n986), .ZN(n778) );
  NAND2_X1 U860 ( .A1(n778), .A2(G868), .ZN(n780) );
  NAND2_X1 U861 ( .A1(n976), .A2(n815), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G123), .A2(n889), .ZN(n781) );
  XNOR2_X1 U864 ( .A(n781), .B(KEYINPUT18), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G135), .A2(n522), .ZN(n782) );
  XOR2_X1 U866 ( .A(KEYINPUT81), .B(n782), .Z(n783) );
  NAND2_X1 U867 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U868 ( .A1(G111), .A2(n888), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G99), .A2(n894), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U871 ( .A1(n788), .A2(n787), .ZN(n937) );
  XNOR2_X1 U872 ( .A(n937), .B(G2096), .ZN(n790) );
  INV_X1 U873 ( .A(G2100), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G156) );
  NAND2_X1 U875 ( .A1(n532), .A2(G93), .ZN(n791) );
  XOR2_X1 U876 ( .A(KEYINPUT83), .B(n791), .Z(n794) );
  NAND2_X1 U877 ( .A1(n792), .A2(G80), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U879 ( .A(KEYINPUT84), .B(n795), .ZN(n801) );
  NAND2_X1 U880 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G55), .A2(n797), .ZN(n798) );
  NAND2_X1 U882 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U883 ( .A1(n801), .A2(n800), .ZN(n814) );
  XOR2_X1 U884 ( .A(n814), .B(KEYINPUT82), .Z(n805) );
  NAND2_X1 U885 ( .A1(G559), .A2(n916), .ZN(n802) );
  XOR2_X1 U886 ( .A(n976), .B(n802), .Z(n812) );
  NAND2_X1 U887 ( .A1(n812), .A2(n803), .ZN(n804) );
  XNOR2_X1 U888 ( .A(n805), .B(n804), .ZN(G145) );
  XNOR2_X1 U889 ( .A(n981), .B(G288), .ZN(n811) );
  XOR2_X1 U890 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n807) );
  XNOR2_X1 U891 ( .A(G166), .B(n814), .ZN(n806) );
  XNOR2_X1 U892 ( .A(n807), .B(n806), .ZN(n808) );
  XOR2_X1 U893 ( .A(n808), .B(G290), .Z(n809) );
  XNOR2_X1 U894 ( .A(G305), .B(n809), .ZN(n810) );
  XNOR2_X1 U895 ( .A(n811), .B(n810), .ZN(n915) );
  XNOR2_X1 U896 ( .A(n812), .B(n915), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U898 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U900 ( .A(KEYINPUT87), .B(n818), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n819) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U905 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U907 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U908 ( .A1(G219), .A2(G220), .ZN(n823) );
  XNOR2_X1 U909 ( .A(KEYINPUT22), .B(n823), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n824), .A2(G96), .ZN(n825) );
  NOR2_X1 U911 ( .A1(G218), .A2(n825), .ZN(n826) );
  XOR2_X1 U912 ( .A(KEYINPUT88), .B(n826), .Z(n838) );
  NAND2_X1 U913 ( .A1(n838), .A2(G2106), .ZN(n830) );
  NAND2_X1 U914 ( .A1(G120), .A2(G108), .ZN(n827) );
  NOR2_X1 U915 ( .A1(G237), .A2(n827), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G69), .A2(n828), .ZN(n837) );
  NAND2_X1 U917 ( .A1(G567), .A2(n837), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n870) );
  NAND2_X1 U919 ( .A1(G483), .A2(G661), .ZN(n831) );
  NOR2_X1 U920 ( .A1(n870), .A2(n831), .ZN(n832) );
  XOR2_X1 U921 ( .A(KEYINPUT89), .B(n832), .Z(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U928 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(G2100), .B(KEYINPUT110), .Z(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT109), .B(G2678), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2072), .Z(n842) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U941 ( .A(KEYINPUT43), .B(G2096), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n848) );
  XOR2_X1 U943 ( .A(G2084), .B(G2078), .Z(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1981), .B(G1971), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(G1976), .B(G1956), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1986), .B(G2474), .Z(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G229) );
  XNOR2_X1 U956 ( .A(G2430), .B(G2454), .ZN(n867) );
  XNOR2_X1 U957 ( .A(KEYINPUT106), .B(G2435), .ZN(n865) );
  XOR2_X1 U958 ( .A(G2451), .B(G2427), .Z(n860) );
  XNOR2_X1 U959 ( .A(G2438), .B(G2446), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n861), .B(G2443), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1341), .B(G1348), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n868), .A2(G14), .ZN(n869) );
  XNOR2_X1 U967 ( .A(KEYINPUT107), .B(n869), .ZN(G401) );
  XOR2_X1 U968 ( .A(KEYINPUT108), .B(n870), .Z(G319) );
  NAND2_X1 U969 ( .A1(G124), .A2(n889), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n871), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G112), .A2(n888), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT112), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G100), .A2(n894), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G136), .A2(n522), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G103), .A2(n894), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G139), .A2(n522), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G115), .A2(n888), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G127), .A2(n889), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT114), .B(n883), .Z(n884) );
  XNOR2_X1 U985 ( .A(KEYINPUT47), .B(n884), .ZN(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n929) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(n937), .ZN(n903) );
  NAND2_X1 U989 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U992 ( .A1(n522), .A2(G142), .ZN(n893) );
  XOR2_X1 U993 ( .A(KEYINPUT113), .B(n893), .Z(n896) );
  NAND2_X1 U994 ( .A1(n894), .A2(G106), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n909) );
  XOR2_X1 U1000 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n929), .B(n910), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n911), .B(G162), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G286), .B(n915), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(G171), .B(n916), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1012 ( .A(n919), .B(n976), .Z(n920) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n920), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n921), .B(KEYINPUT49), .ZN(n925) );
  INV_X1 U1016 ( .A(G401), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n922), .A2(G319), .ZN(n923) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(n923), .Z(n924) );
  NOR2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(n981), .ZN(G299) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n928) );
  XNOR2_X1 U1026 ( .A(KEYINPUT120), .B(n928), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G2072), .B(n929), .Z(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT50), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n950) );
  XNOR2_X1 U1031 ( .A(G2084), .B(G160), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT119), .B(n935), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n941) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n946) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT51), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n972) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n972), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n966) );
  XOR2_X1 U1047 ( .A(G1991), .B(G25), .Z(n954) );
  NAND2_X1 U1048 ( .A1(n954), .A2(G28), .ZN(n963) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(KEYINPUT121), .B(n967), .Z(n970) );
  XOR2_X1 U1060 ( .A(KEYINPUT54), .B(G34), .Z(n968) );
  XNOR2_X1 U1061 ( .A(G2084), .B(n968), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n972), .B(n971), .ZN(n974) );
  INV_X1 U1064 ( .A(G29), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n975), .ZN(n1028) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1068 ( .A(G301), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(n976), .B(G1341), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n998) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n981), .B(G1956), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n996) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1081 ( .A(KEYINPUT122), .B(n993), .Z(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT57), .B(n994), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  INV_X1 U1086 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .Z(n1001) );
  XNOR2_X1 U1088 ( .A(G4), .B(n1001), .ZN(n1008) );
  XOR2_X1 U1089 ( .A(G1341), .B(G19), .Z(n1005) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT123), .B(n1006), .Z(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1009), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1971), .B(KEYINPUT124), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G22), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1114 ( .A(n1031), .B(KEYINPUT62), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(KEYINPUT125), .B(n1032), .ZN(G311) );
  XOR2_X1 U1116 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

