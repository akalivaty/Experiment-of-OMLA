

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X2 U321 ( .A1(n520), .A2(n414), .ZN(n569) );
  INV_X1 U322 ( .A(n531), .ZN(n412) );
  XOR2_X1 U323 ( .A(n574), .B(KEYINPUT41), .Z(n563) );
  NAND2_X1 U324 ( .A1(n412), .A2(n522), .ZN(n413) );
  XNOR2_X1 U325 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U326 ( .A(n413), .B(KEYINPUT54), .ZN(n414) );
  XNOR2_X1 U327 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U328 ( .A(KEYINPUT98), .B(n471), .Z(n520) );
  XNOR2_X1 U329 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XNOR2_X1 U330 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT97), .B(KEYINPUT92), .Z(n290) );
  XNOR2_X1 U332 ( .A(G162GAT), .B(KEYINPUT95), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G57GAT), .Z(n320) );
  XOR2_X1 U335 ( .A(n291), .B(n320), .Z(n297) );
  XOR2_X1 U336 ( .A(G113GAT), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U337 ( .A(G29GAT), .B(G134GAT), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n292), .B(G85GAT), .ZN(n346) );
  XOR2_X1 U339 ( .A(KEYINPUT0), .B(G127GAT), .Z(n446) );
  XOR2_X1 U340 ( .A(n346), .B(n446), .Z(n294) );
  NAND2_X1 U341 ( .A1(G225GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n387), .B(n295), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U345 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n299) );
  XNOR2_X1 U346 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n301), .B(n300), .Z(n310) );
  XNOR2_X1 U349 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n302), .B(KEYINPUT89), .ZN(n303) );
  XOR2_X1 U351 ( .A(n303), .B(KEYINPUT2), .Z(n305) );
  XNOR2_X1 U352 ( .A(G141GAT), .B(G148GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n422) );
  XOR2_X1 U354 ( .A(KEYINPUT4), .B(KEYINPUT96), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n422), .B(n308), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n471) );
  XOR2_X1 U359 ( .A(G99GAT), .B(G106GAT), .Z(n330) );
  XOR2_X1 U360 ( .A(G71GAT), .B(KEYINPUT13), .Z(n362) );
  XOR2_X1 U361 ( .A(n330), .B(n362), .Z(n312) );
  NAND2_X1 U362 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U364 ( .A(KEYINPUT70), .B(KEYINPUT73), .Z(n314) );
  XNOR2_X1 U365 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(n316), .B(n315), .Z(n322) );
  XOR2_X1 U368 ( .A(G92GAT), .B(G85GAT), .Z(n318) );
  XNOR2_X1 U369 ( .A(G148GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U373 ( .A(n323), .B(KEYINPUT72), .Z(n327) );
  XOR2_X1 U374 ( .A(G64GAT), .B(KEYINPUT71), .Z(n325) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G204GAT), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n408) );
  XNOR2_X1 U377 ( .A(n408), .B(KEYINPUT32), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n574) );
  XNOR2_X1 U379 ( .A(G92GAT), .B(G218GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n332) );
  INV_X1 U382 ( .A(n332), .ZN(n404) );
  NAND2_X1 U383 ( .A1(n330), .A2(n404), .ZN(n334) );
  INV_X1 U384 ( .A(n330), .ZN(n331) );
  NAND2_X1 U385 ( .A1(n332), .A2(n331), .ZN(n333) );
  NAND2_X1 U386 ( .A1(n334), .A2(n333), .ZN(n336) );
  AND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U390 ( .A(n418), .B(KEYINPUT65), .ZN(n338) );
  INV_X1 U391 ( .A(KEYINPUT11), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT74), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U395 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n345), .B(KEYINPUT7), .ZN(n388) );
  XNOR2_X1 U398 ( .A(n388), .B(n346), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n558) );
  XNOR2_X1 U400 ( .A(KEYINPUT75), .B(n558), .ZN(n544) );
  XNOR2_X1 U401 ( .A(n544), .B(KEYINPUT36), .ZN(n580) );
  XOR2_X1 U402 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n350) );
  XNOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT77), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n370) );
  XOR2_X1 U405 ( .A(G64GAT), .B(G57GAT), .Z(n352) );
  XNOR2_X1 U406 ( .A(G1GAT), .B(G211GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(KEYINPUT76), .Z(n354) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(KEYINPUT82), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U411 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U412 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n358) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT81), .B(n359), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U417 ( .A(G22GAT), .B(G78GAT), .Z(n426) );
  XOR2_X1 U418 ( .A(n362), .B(n426), .Z(n364) );
  XNOR2_X1 U419 ( .A(G183GAT), .B(G155GAT), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U421 ( .A(n366), .B(n365), .Z(n368) );
  XNOR2_X1 U422 ( .A(G15GAT), .B(G127GAT), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U424 ( .A(n370), .B(n369), .Z(n489) );
  NAND2_X1 U425 ( .A1(n580), .A2(n489), .ZN(n372) );
  XOR2_X1 U426 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n373) );
  NAND2_X1 U428 ( .A1(n574), .A2(n373), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n374), .B(KEYINPUT119), .ZN(n391) );
  XOR2_X1 U430 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n376) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U433 ( .A(n377), .B(KEYINPUT69), .Z(n385) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G50GAT), .Z(n379) );
  XNOR2_X1 U435 ( .A(G29GAT), .B(G36GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U437 ( .A(KEYINPUT68), .B(G197GAT), .Z(n381) );
  XNOR2_X1 U438 ( .A(G141GAT), .B(G22GAT), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XOR2_X1 U443 ( .A(n386), .B(n401), .Z(n390) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n570) );
  NAND2_X1 U446 ( .A1(n391), .A2(n570), .ZN(n398) );
  XOR2_X1 U447 ( .A(KEYINPUT118), .B(KEYINPUT47), .Z(n396) );
  NOR2_X1 U448 ( .A1(n570), .A2(n563), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n392), .B(KEYINPUT46), .ZN(n393) );
  NOR2_X1 U450 ( .A1(n489), .A2(n393), .ZN(n394) );
  NAND2_X1 U451 ( .A1(n394), .A2(n558), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U453 ( .A1(n398), .A2(n397), .ZN(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT48), .B(n399), .Z(n531) );
  XOR2_X1 U455 ( .A(G197GAT), .B(KEYINPUT21), .Z(n400) );
  XOR2_X1 U456 ( .A(G211GAT), .B(n400), .Z(n417) );
  XOR2_X1 U457 ( .A(KEYINPUT99), .B(n401), .Z(n403) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U460 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U461 ( .A(G183GAT), .B(KEYINPUT17), .Z(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n434) );
  XNOR2_X1 U464 ( .A(n434), .B(n408), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n417), .B(n411), .ZN(n522) );
  INV_X1 U467 ( .A(n522), .ZN(n458) );
  XOR2_X1 U468 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U469 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n432) );
  XOR2_X1 U471 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n430) );
  XOR2_X1 U475 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n424) );
  XNOR2_X1 U476 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U478 ( .A(n425), .B(G106GAT), .Z(n428) );
  XNOR2_X1 U479 ( .A(n426), .B(G218GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n432), .B(n431), .ZN(n464) );
  NAND2_X1 U483 ( .A1(n569), .A2(n464), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n433), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U485 ( .A(G169GAT), .B(n434), .Z(n436) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n452) );
  XOR2_X1 U488 ( .A(G71GAT), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U489 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U491 ( .A(G120GAT), .B(KEYINPUT83), .Z(n440) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(G113GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT64), .Z(n444) );
  XNOR2_X1 U496 ( .A(G99GAT), .B(G190GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n445), .B(G134GAT), .Z(n448) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n525) );
  NAND2_X1 U503 ( .A1(n453), .A2(n525), .ZN(n566) );
  INV_X1 U504 ( .A(n566), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n454), .A2(n544), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT105), .B(KEYINPUT34), .Z(n478) );
  INV_X1 U507 ( .A(n570), .ZN(n505) );
  NAND2_X1 U508 ( .A1(n574), .A2(n505), .ZN(n492) );
  INV_X1 U509 ( .A(n489), .ZN(n577) );
  NOR2_X1 U510 ( .A1(n544), .A2(n577), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT16), .ZN(n475) );
  INV_X1 U512 ( .A(n525), .ZN(n533) );
  XOR2_X1 U513 ( .A(n458), .B(KEYINPUT27), .Z(n467) );
  NAND2_X1 U514 ( .A1(n520), .A2(n467), .ZN(n530) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n464), .Z(n532) );
  NOR2_X1 U516 ( .A1(n530), .A2(n532), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n533), .A2(n459), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT100), .ZN(n474) );
  NAND2_X1 U519 ( .A1(n525), .A2(n522), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n461), .A2(n464), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT102), .ZN(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .Z(n469) );
  NOR2_X1 U523 ( .A1(n525), .A2(n464), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT26), .B(n465), .Z(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT101), .B(n466), .ZN(n568) );
  NAND2_X1 U526 ( .A1(n467), .A2(n568), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT103), .B(n470), .Z(n472) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n487) );
  NAND2_X1 U531 ( .A1(n475), .A2(n487), .ZN(n506) );
  NOR2_X1 U532 ( .A1(n492), .A2(n506), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT104), .B(n476), .ZN(n484) );
  NAND2_X1 U534 ( .A1(n520), .A2(n484), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n484), .A2(n522), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT106), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U541 ( .A1(n484), .A2(n525), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  XOR2_X1 U543 ( .A(G22GAT), .B(KEYINPUT107), .Z(n486) );
  NAND2_X1 U544 ( .A1(n484), .A2(n532), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  NAND2_X1 U546 ( .A1(n580), .A2(n487), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(KEYINPUT108), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n519) );
  NOR2_X1 U550 ( .A1(n492), .A2(n519), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(KEYINPUT38), .ZN(n502) );
  NAND2_X1 U552 ( .A1(n520), .A2(n502), .ZN(n495) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n497) );
  NAND2_X1 U556 ( .A1(n502), .A2(n522), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n500) );
  NAND2_X1 U560 ( .A1(n502), .A2(n525), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n532), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT112), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT113), .Z(n508) );
  OR2_X1 U567 ( .A1(n505), .A2(n563), .ZN(n518) );
  NOR2_X1 U568 ( .A1(n506), .A2(n518), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n513), .A2(n520), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n522), .A2(n513), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n525), .A2(n513), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT114), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT115), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U578 ( .A1(n513), .A2(n532), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT116), .Z(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n520), .A2(n527), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT117), .Z(n524) );
  NAND2_X1 U586 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n527), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n548) );
  NOR2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n548), .A2(n534), .ZN(n543) );
  NOR2_X1 U596 ( .A1(n570), .A2(n543), .ZN(n536) );
  XNOR2_X1 U597 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  NOR2_X1 U600 ( .A1(n563), .A2(n543), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n577), .A2(n543), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT122), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  INV_X1 U608 ( .A(n543), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n568), .ZN(n557) );
  NOR2_X1 U612 ( .A1(n570), .A2(n557), .ZN(n550) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT123), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT124), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n554) );
  NOR2_X1 U618 ( .A1(n563), .A2(n557), .ZN(n553) );
  XOR2_X1 U619 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n577), .A2(n557), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT125), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n559), .Z(G1347GAT) );
  NOR2_X1 U625 ( .A1(n570), .A2(n566), .ZN(n560) );
  XOR2_X1 U626 ( .A(G169GAT), .B(n560), .Z(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT126), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n565) );
  NOR2_X1 U630 ( .A1(n563), .A2(n566), .ZN(n564) );
  XOR2_X1 U631 ( .A(n565), .B(n564), .Z(G1349GAT) );
  NOR2_X1 U632 ( .A1(n577), .A2(n566), .ZN(n567) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n579) );
  NOR2_X1 U635 ( .A1(n570), .A2(n579), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n583) );
  INV_X1 U645 ( .A(n579), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

