//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n212), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G50), .B2(G226), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n209), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n225), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(G20), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT7), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  AOI211_X1 g0055(.A(new_n255), .B(G20), .C1(new_n250), .C2(new_n252), .ZN(new_n256));
  OAI21_X1  g0056(.A(G68), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  INV_X1    g0058(.A(G68), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n260), .B2(new_n202), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G159), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n248), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT71), .B1(new_n253), .B2(KEYINPUT7), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n255), .C1(new_n271), .C2(G20), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n256), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT16), .B(new_n265), .C1(new_n273), .C2(new_n259), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n247), .B1(new_n275), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n278), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n268), .A2(new_n274), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n249), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  OR2_X1    g0091(.A1(G223), .A2(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n271), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G87), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G232), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n295), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NOR4_X1   g0106(.A1(new_n295), .A2(new_n299), .A3(new_n302), .A4(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT18), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n287), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n255), .B1(new_n271), .B2(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n250), .A2(new_n252), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n259), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n267), .B1(new_n314), .B2(new_n264), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n274), .A2(new_n247), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n285), .A2(new_n286), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n305), .A2(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT18), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n293), .A2(new_n294), .ZN(new_n322));
  INV_X1    g0122(.A(new_n289), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  INV_X1    g0125(.A(new_n299), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n301), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n303), .B2(G200), .ZN(new_n328));
  INV_X1    g0128(.A(new_n274), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n315), .A2(new_n247), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n317), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT17), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT73), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n316), .A2(new_n337), .A3(new_n317), .A4(new_n328), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT74), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n287), .A2(new_n340), .A3(new_n337), .A4(new_n328), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n321), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n301), .B1(new_n297), .B2(new_n221), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G238), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n271), .B(new_n346), .C1(new_n298), .C2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n323), .C1(G107), .C2(new_n271), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n325), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n345), .B2(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n276), .A2(G77), .ZN(new_n353));
  XOR2_X1   g0153(.A(new_n353), .B(KEYINPUT69), .Z(new_n354));
  INV_X1    g0154(.A(new_n281), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n220), .ZN(new_n356));
  INV_X1    g0156(.A(new_n262), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n226), .A2(G33), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n280), .A2(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n226), .A2(new_n220), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n247), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n354), .A2(new_n356), .A3(new_n363), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n350), .A2(new_n352), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n343), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n281), .A2(G50), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT67), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n262), .A2(G150), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT67), .B(G20), .C1(new_n201), .C2(new_n203), .ZN(new_n372));
  INV_X1    g0172(.A(new_n360), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n278), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n370), .A2(new_n371), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n367), .B1(new_n375), .B2(new_n247), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n276), .A2(G50), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT9), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n301), .B1(new_n297), .B2(new_n290), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT66), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G222), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G223), .A2(G1698), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n271), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n323), .C1(G77), .C2(new_n271), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n301), .B(KEYINPUT66), .C1(new_n297), .C2(new_n290), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(new_n325), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(G200), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT70), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT70), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n394), .A3(G200), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n379), .A2(new_n380), .A3(new_n391), .A4(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n378), .A2(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT9), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n376), .B2(new_n377), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n391), .B(new_n396), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n390), .A2(new_n304), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n378), .B(new_n404), .C1(G179), .C2(new_n390), .ZN(new_n405));
  INV_X1    g0205(.A(G50), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n357), .A2(new_n406), .B1(new_n360), .B2(new_n220), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n226), .A2(G68), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n247), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT11), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n276), .A2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n275), .A3(G13), .ZN(new_n414));
  XOR2_X1   g0214(.A(new_n414), .B(KEYINPUT12), .Z(new_n415));
  NOR3_X1   g0215(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(G226), .A2(G1698), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n298), .B2(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n271), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n323), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n289), .A2(G238), .A3(new_n296), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n301), .A4(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n418), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n301), .B(new_n424), .C1(new_n426), .C2(new_n289), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n416), .B1(new_n429), .B2(new_n325), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n351), .B1(new_n425), .B2(new_n428), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n429), .B2(G169), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n429), .A2(new_n306), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n429), .A2(new_n433), .A3(G169), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n416), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n349), .A2(new_n304), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n345), .A2(new_n306), .A3(new_n348), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n364), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n403), .A2(new_n405), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n366), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n281), .A2(G116), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n249), .A2(G1), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n225), .B(new_n246), .C1(new_n448), .C2(KEYINPUT75), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n275), .A2(KEYINPUT75), .A3(G33), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n281), .A2(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n226), .C1(G33), .C2(new_n214), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT81), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(new_n249), .B2(G97), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n458), .A3(new_n454), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n450), .A2(G20), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n459), .A3(new_n460), .A4(new_n247), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n455), .A2(KEYINPUT81), .B1(new_n225), .B2(new_n246), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n460), .A4(new_n459), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n447), .B(new_n453), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n275), .B(G45), .C1(new_n288), .C2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT5), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT77), .B1(new_n469), .B2(G41), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT77), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n288), .A3(KEYINPUT5), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT78), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT78), .B1(new_n470), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g0274(.A(G274), .B(new_n468), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G264), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n271), .B(new_n476), .C1(new_n215), .C2(G1698), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n312), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n323), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(new_n472), .ZN(new_n481));
  OAI211_X1 g0281(.A(G270), .B(new_n289), .C1(new_n481), .C2(new_n467), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n466), .A2(new_n306), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n483), .A2(new_n325), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(G200), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n466), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(G169), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n466), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n489), .B(KEYINPUT21), .C1(new_n466), .C2(new_n490), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n484), .B(new_n488), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n250), .A2(new_n252), .A3(G244), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(new_n250), .A3(new_n252), .A4(G244), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n454), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n250), .A2(new_n252), .A3(G250), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n384), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n323), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n470), .A2(new_n472), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n323), .B1(new_n505), .B2(new_n468), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G257), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n475), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n355), .A2(new_n214), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT76), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n449), .B2(new_n452), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT75), .B1(new_n275), .B2(G33), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n247), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(KEYINPUT76), .A3(new_n281), .A4(new_n451), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n512), .A2(new_n515), .A3(G97), .ZN(new_n516));
  OAI21_X1  g0316(.A(G107), .B1(new_n254), .B2(new_n256), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n214), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n226), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n262), .A2(G77), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n516), .B1(new_n527), .B2(new_n247), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n504), .A2(G190), .A3(new_n475), .A4(new_n507), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n509), .A2(new_n510), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n512), .A2(new_n515), .A3(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n519), .B1(new_n311), .B2(new_n313), .ZN(new_n532));
  INV_X1    g0332(.A(new_n526), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n532), .A2(new_n533), .A3(new_n524), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n510), .B(new_n531), .C1(new_n534), .C2(new_n248), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n508), .A2(new_n304), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n504), .A2(new_n306), .A3(new_n475), .A4(new_n507), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n530), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n355), .B(new_n519), .C1(KEYINPUT85), .C2(KEYINPUT25), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n512), .A2(new_n515), .A3(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT23), .B1(new_n519), .B2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n519), .A2(KEYINPUT23), .A3(G20), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(new_n373), .B2(G116), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n250), .A2(new_n252), .A3(new_n226), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(G87), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n250), .A2(new_n252), .A3(new_n226), .A4(G87), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT84), .B1(new_n554), .B2(KEYINPUT83), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n552), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n548), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT24), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n548), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n544), .B1(new_n562), .B2(new_n247), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n213), .A2(new_n384), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n215), .A2(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n250), .A2(new_n564), .A3(new_n252), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n249), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n506), .A2(G264), .B1(new_n568), .B2(new_n323), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n475), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n351), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G190), .B2(new_n570), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n539), .B1(new_n563), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G45), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n213), .B1(new_n574), .B2(G1), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n275), .A2(new_n300), .A3(G45), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n289), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n221), .A2(G1698), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n250), .A2(new_n578), .A3(new_n252), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G116), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n577), .B1(new_n582), .B2(new_n289), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n325), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n212), .A2(new_n214), .A3(new_n519), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n420), .A2(new_n226), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT19), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n360), .B2(new_n214), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n271), .A2(new_n226), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n588), .B(new_n590), .C1(new_n591), .C2(new_n259), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n247), .B1(new_n355), .B2(new_n359), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n512), .A2(new_n515), .A3(G87), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n583), .A2(G200), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n289), .B1(new_n580), .B2(new_n581), .ZN(new_n597));
  INV_X1    g0397(.A(new_n577), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n585), .A2(new_n595), .A3(new_n596), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n599), .A2(new_n304), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n597), .A2(new_n598), .A3(new_n306), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT79), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n583), .A2(G169), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT79), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(G179), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n512), .A2(new_n515), .A3(new_n358), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n593), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n603), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n562), .A2(new_n247), .ZN(new_n615));
  INV_X1    g0415(.A(new_n544), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT86), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n569), .A2(new_n618), .A3(G179), .A4(new_n475), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT86), .B1(new_n570), .B2(G169), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n570), .A2(new_n306), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n446), .A2(new_n495), .A3(new_n573), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT87), .ZN(G372));
  AOI21_X1  g0425(.A(new_n484), .B1(new_n493), .B2(new_n494), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n248), .B1(new_n559), .B2(new_n561), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n627), .B2(new_n544), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n607), .A2(new_n609), .B1(new_n593), .B2(new_n611), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT88), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT88), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n593), .A2(new_n596), .A3(new_n594), .A4(new_n600), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n629), .A2(new_n573), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n603), .A2(new_n613), .ZN(new_n639));
  INV_X1    g0439(.A(new_n538), .ZN(new_n640));
  XNOR2_X1  g0440(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n538), .B1(new_n633), .B2(new_n636), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n638), .A2(new_n631), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n446), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n439), .A2(new_n440), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n432), .B2(new_n444), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT73), .B1(new_n331), .B2(KEYINPUT17), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n331), .A2(KEYINPUT73), .A3(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n342), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n321), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n403), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n405), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(G13), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G20), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n275), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT90), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n495), .B1(new_n466), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n667), .A2(new_n466), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n626), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n617), .B1(new_n622), .B2(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n563), .A2(new_n572), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n628), .B2(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n617), .A2(new_n622), .A3(new_n667), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n626), .A2(new_n666), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n679), .A2(new_n673), .A3(new_n674), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n207), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n586), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n228), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n640), .ZN(new_n689));
  INV_X1    g0489(.A(new_n641), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n614), .B2(new_n538), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n638), .A2(new_n692), .A3(new_n631), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n667), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n645), .A2(new_n696), .A3(new_n667), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n623), .A2(new_n495), .A3(new_n573), .A4(new_n667), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT31), .ZN(new_n701));
  INV_X1    g0501(.A(new_n508), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n609), .A2(new_n483), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(KEYINPUT30), .A4(new_n569), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n569), .A2(new_n504), .A3(new_n475), .A4(new_n507), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n605), .A2(new_n480), .A3(new_n482), .A4(new_n475), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT91), .B1(new_n508), .B2(new_n570), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n508), .A2(new_n570), .A3(KEYINPUT91), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n599), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n483), .A2(new_n306), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT92), .B(new_n701), .C1(new_n715), .C2(new_n667), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n704), .A2(new_n708), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n570), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n583), .B(new_n714), .C1(new_n718), .C2(new_n710), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n667), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n720), .B2(KEYINPUT31), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n700), .A2(new_n716), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n699), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n688), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR3_X1   g0528(.A1(new_n657), .A2(new_n574), .A3(G20), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n683), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n672), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n670), .ZN(new_n735));
  INV_X1    g0535(.A(new_n733), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n225), .B1(G20), .B2(new_n304), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n226), .A2(new_n306), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n351), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n325), .A3(new_n351), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G326), .A2(new_n741), .B1(new_n743), .B2(G311), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n325), .A3(G200), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT33), .B(G317), .Z(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n226), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n271), .B1(new_n751), .B2(G329), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n351), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n740), .A2(G200), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n747), .B(new_n759), .C1(G322), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n226), .B1(new_n749), .B2(G190), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT95), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT95), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n753), .A2(G20), .A3(G190), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n761), .B1(new_n567), .B2(new_n765), .C1(new_n478), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n760), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n770), .A2(new_n258), .B1(new_n259), .B2(new_n745), .ZN(new_n771));
  INV_X1    g0571(.A(new_n757), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n769), .B(new_n771), .C1(G107), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT32), .B1(new_n750), .B2(new_n768), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n766), .A2(new_n212), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n312), .ZN(new_n776));
  INV_X1    g0576(.A(new_n741), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n777), .A2(new_n406), .B1(new_n220), .B2(new_n742), .ZN(new_n778));
  INV_X1    g0578(.A(new_n765), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(G97), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n773), .A2(new_n774), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n738), .B1(new_n767), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n737), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n682), .A2(new_n271), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n229), .A2(new_n574), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n241), .C2(new_n574), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n271), .A2(new_n207), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G116), .B2(new_n207), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n782), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n785), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n670), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n735), .B1(new_n736), .B2(new_n795), .ZN(G396));
  NAND2_X1  g0596(.A1(new_n645), .A2(new_n667), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n666), .A2(new_n364), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n365), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n444), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n444), .A2(new_n666), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n797), .B(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(new_n725), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n736), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n757), .A2(new_n212), .B1(new_n519), .B2(new_n766), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n742), .A2(new_n450), .B1(new_n745), .B2(new_n758), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n770), .A2(new_n567), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n312), .B1(new_n750), .B2(new_n811), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n813), .B1(new_n214), .B2(new_n765), .C1(new_n478), .C2(new_n777), .ZN(new_n814));
  INV_X1    g0614(.A(new_n745), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n760), .B1(new_n815), .B2(G150), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n741), .A2(G137), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n768), .C2(new_n742), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n271), .B1(new_n406), .B2(new_n766), .C1(new_n765), .C2(new_n258), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n819), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n772), .A2(G68), .B1(G132), .B2(new_n751), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n738), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n737), .A2(new_n783), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT96), .Z(new_n828));
  AOI21_X1  g0628(.A(new_n826), .B1(new_n220), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n733), .B(new_n829), .C1(new_n804), .C2(new_n784), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n807), .A2(new_n830), .ZN(G384));
  INV_X1    g0631(.A(KEYINPUT99), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n287), .B2(new_n664), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n318), .A2(KEYINPUT99), .A3(new_n663), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n318), .A2(new_n319), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n331), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n265), .B1(new_n273), .B2(new_n259), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n267), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n247), .A3(new_n274), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n841), .A2(new_n283), .B1(new_n308), .B2(new_n664), .ZN(new_n842));
  INV_X1    g0642(.A(new_n331), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n310), .A2(new_n320), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n651), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n664), .B1(new_n841), .B2(new_n283), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT98), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT98), .ZN(new_n850));
  INV_X1    g0650(.A(new_n848), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(new_n651), .C2(new_n846), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n845), .B(KEYINPUT38), .C1(new_n849), .C2(new_n852), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  INV_X1    g0658(.A(new_n845), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n850), .B1(new_n343), .B2(new_n851), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n334), .A2(new_n335), .B1(new_n339), .B2(new_n341), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT98), .B(new_n848), .C1(new_n861), .C2(new_n321), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n854), .B(new_n859), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n847), .A2(new_n833), .A3(new_n834), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n835), .A2(new_n837), .A3(new_n331), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n838), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n647), .A2(new_n666), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n857), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n846), .A2(new_n663), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n855), .A2(new_n856), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n802), .B1(new_n797), .B2(new_n803), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n440), .B(new_n666), .C1(new_n439), .C2(new_n432), .ZN(new_n875));
  INV_X1    g0675(.A(new_n432), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n666), .A2(new_n440), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT14), .B(new_n304), .C1(new_n425), .C2(new_n428), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n434), .A2(new_n878), .A3(new_n436), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n876), .B(new_n877), .C1(new_n879), .C2(new_n416), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n872), .B1(new_n873), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT100), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n871), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n871), .B2(new_n884), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n645), .A2(new_n696), .A3(new_n667), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n696), .B1(new_n693), .B2(new_n667), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n446), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(new_n446), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n655), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n888), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n720), .B(new_n701), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n803), .B(new_n881), .C1(new_n898), .C2(new_n700), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n860), .A2(new_n862), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n900), .B2(new_n845), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n901), .B2(new_n863), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n864), .A2(new_n867), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n854), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n856), .A2(new_n905), .B1(new_n899), .B2(KEYINPUT102), .ZN(new_n906));
  INV_X1    g0706(.A(new_n700), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n701), .B1(new_n715), .B2(new_n667), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n721), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n804), .B(new_n882), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n903), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n902), .A2(new_n903), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n898), .A2(new_n700), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n446), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(G330), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n897), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n275), .B2(new_n658), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n228), .A2(new_n220), .A3(new_n260), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n201), .A2(new_n259), .ZN(new_n921));
  OAI211_X1 g0721(.A(G1), .B(new_n657), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n522), .A2(new_n523), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n450), .B1(new_n923), .B2(KEYINPUT35), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(new_n227), .C1(KEYINPUT35), .C2(new_n923), .ZN(new_n925));
  XOR2_X1   g0725(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n919), .A2(new_n922), .A3(new_n927), .ZN(G367));
  OR2_X1    g0728(.A1(new_n667), .A2(new_n595), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n631), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n637), .B2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT43), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n666), .A2(new_n535), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n538), .A3(new_n530), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n680), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n538), .B1(new_n936), .B2(new_n628), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n667), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n934), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n932), .B2(new_n931), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(new_n934), .A3(new_n940), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT103), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n640), .A2(new_n666), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n936), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n677), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n947), .A2(new_n952), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n683), .B(new_n955), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n680), .A2(new_n678), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n950), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n950), .C1(KEYINPUT106), .C2(KEYINPUT44), .ZN(new_n962));
  AND2_X1   g0762(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n677), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n680), .B1(new_n676), .B2(new_n679), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n671), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n726), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n957), .B1(new_n973), .B2(new_n727), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n953), .B(new_n954), .C1(new_n974), .C2(new_n732), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n757), .A2(new_n214), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n271), .B(new_n976), .C1(G317), .C2(new_n751), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT107), .Z(new_n978));
  OAI22_X1  g0778(.A1(new_n770), .A2(new_n478), .B1(new_n567), .B2(new_n745), .ZN(new_n979));
  INV_X1    g0779(.A(new_n766), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G116), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT46), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n981), .A2(new_n982), .B1(G283), .B2(new_n743), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n811), .B2(new_n777), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n979), .B(new_n984), .C1(G107), .C2(new_n779), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n978), .B(new_n985), .C1(new_n982), .C2(new_n981), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n772), .A2(G77), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G143), .A2(new_n741), .B1(new_n815), .B2(G159), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n312), .B1(new_n751), .B2(G137), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n980), .A2(G58), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT108), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n779), .A2(G68), .ZN(new_n993));
  INV_X1    g0793(.A(G150), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n770), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n991), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n201), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n996), .B1(new_n992), .B2(new_n995), .C1(new_n997), .C2(new_n742), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n986), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT109), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n736), .B1(new_n1001), .B2(new_n737), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n787), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n786), .B1(new_n207), .B2(new_n359), .C1(new_n237), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n931), .A2(new_n785), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n975), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT110), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n975), .A2(KEYINPUT110), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(G387));
  AOI22_X1  g0811(.A1(G317), .A2(new_n760), .B1(new_n815), .B2(G311), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n741), .A2(G322), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n478), .C2(new_n742), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(new_n1016), .B1(G283), .B2(new_n779), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n567), .B2(new_n766), .C1(new_n1016), .C2(new_n1015), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT49), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n751), .A2(G326), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n271), .B1(new_n772), .B2(G116), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n760), .B1(new_n743), .B2(G68), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n768), .B2(new_n777), .C1(new_n280), .C2(new_n745), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT112), .B(G150), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n976), .B(new_n1026), .C1(new_n751), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n980), .A2(G77), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n779), .A2(new_n358), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1024), .B1(new_n312), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n278), .A2(new_n406), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT50), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n685), .A2(KEYINPUT111), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n574), .B1(new_n685), .B2(KEYINPUT111), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n787), .C1(new_n234), .C2(new_n574), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(G107), .B2(new_n207), .C1(new_n685), .C2(new_n791), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1032), .A2(new_n737), .B1(new_n786), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n733), .C1(new_n676), .C2(new_n794), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n732), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n971), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n683), .B1(new_n727), .B2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1042), .B1(new_n1043), .B2(new_n971), .C1(new_n1045), .C2(new_n972), .ZN(G393));
  NAND2_X1  g0846(.A1(new_n968), .A2(new_n969), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n972), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n684), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1049), .A2(new_n973), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n786), .B1(new_n214), .B2(new_n207), .C1(new_n244), .C2(new_n1003), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n280), .A2(new_n742), .B1(new_n997), .B2(new_n745), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n271), .B1(new_n766), .B2(new_n259), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n772), .C2(G87), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n779), .A2(G77), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n751), .A2(G143), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G150), .A2(new_n741), .B1(new_n760), .B2(G159), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n742), .A2(new_n567), .B1(new_n745), .B2(new_n478), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n312), .B1(new_n766), .B2(new_n758), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n772), .C2(G107), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n751), .A2(G322), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n741), .A2(G317), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n770), .B2(new_n811), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT52), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n779), .B2(G116), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1057), .A2(new_n1059), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n736), .B1(new_n1070), .B2(new_n737), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1051), .B(new_n1071), .C1(new_n949), .C2(new_n794), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1047), .B2(new_n1043), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1050), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NAND4_X1  g0875(.A1(new_n724), .A2(G330), .A3(new_n804), .A4(new_n882), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n856), .A2(new_n905), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n693), .A2(new_n667), .A3(new_n800), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n802), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n882), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n870), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT39), .B1(new_n856), .B2(new_n905), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n901), .A2(new_n863), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(KEYINPUT39), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n870), .B1(new_n874), .B2(new_n882), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1076), .B(new_n1082), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n803), .B1(new_n898), .B2(new_n700), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(G330), .A3(new_n882), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n857), .B2(new_n869), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1082), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1087), .A2(new_n1093), .A3(new_n732), .ZN(new_n1094));
  INV_X1    g0894(.A(G132), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n271), .B1(new_n770), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n980), .A2(new_n1027), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(new_n201), .C2(new_n772), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n815), .A2(G137), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n751), .A2(G125), .ZN(new_n1101));
  INV_X1    g0901(.A(G128), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n777), .A2(new_n1102), .B1(new_n742), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G159), .B2(new_n779), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1055), .B1(new_n450), .B2(new_n770), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G283), .A2(new_n741), .B1(new_n815), .B2(G107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n214), .B2(new_n742), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G68), .B2(new_n772), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n271), .B(new_n775), .C1(G294), .C2(new_n751), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n738), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n280), .B2(new_n828), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n733), .B(new_n1116), .C1(new_n1085), .C2(new_n784), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1094), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n446), .A2(G330), .A3(new_n914), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT114), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT114), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n446), .A2(new_n1122), .A3(new_n914), .A4(G330), .ZN(new_n1123));
  AOI221_X4 g0923(.A(new_n654), .B1(new_n1121), .B2(new_n1123), .C1(new_n892), .C2(new_n894), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1088), .A2(G330), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n881), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1079), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1076), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n874), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n724), .A2(G330), .A3(new_n804), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n899), .A2(G330), .B1(new_n1130), .B2(new_n881), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1128), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AOI221_X4 g0932(.A(KEYINPUT115), .B1(new_n1124), .B2(new_n1132), .C1(new_n1087), .C2(new_n1093), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT115), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1087), .A2(new_n1093), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n655), .A3(new_n895), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n893), .B1(new_n698), .B2(new_n446), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n894), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n655), .B(new_n1136), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1076), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n882), .B1(new_n1088), .B2(G330), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1130), .A2(new_n881), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1089), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1145), .A2(new_n1127), .B1(new_n1147), .B2(new_n874), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n1087), .A3(new_n1093), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1150), .A2(new_n683), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT116), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n901), .A2(new_n863), .A3(new_n858), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1153), .A2(new_n1083), .B1(new_n870), .B2(new_n883), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1089), .B1(new_n1154), .B2(new_n1082), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1091), .A2(new_n1143), .A3(new_n1092), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1137), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(KEYINPUT115), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1135), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1159));
  AND4_X1   g0959(.A1(KEYINPUT116), .A2(new_n1151), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1119), .B1(new_n1152), .B2(new_n1160), .ZN(G378));
  NAND3_X1  g0961(.A1(new_n871), .A2(new_n884), .A3(new_n885), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n871), .A2(new_n884), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT100), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT122), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n403), .A2(new_n1165), .A3(new_n405), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n403), .B2(new_n405), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n378), .A2(new_n663), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n913), .B2(G330), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1088), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1077), .A2(new_n912), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n910), .B1(new_n855), .B2(new_n856), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(G330), .C1(new_n1179), .C2(KEYINPUT40), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1174), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1173), .B(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1162), .B(new_n1164), .C1(new_n1176), .C2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n913), .A2(G330), .A3(new_n1175), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n886), .C2(new_n887), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n888), .B(KEYINPUT123), .C1(new_n1183), .C2(new_n1176), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1150), .A2(new_n1124), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1184), .A2(new_n1188), .B1(new_n1124), .B2(new_n1150), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n684), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1189), .A2(new_n732), .A3(new_n1190), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n751), .A2(G283), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1029), .A2(new_n1199), .A3(new_n288), .A4(new_n312), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G107), .A2(new_n760), .B1(new_n815), .B2(G97), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n450), .B2(new_n777), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(new_n358), .C2(new_n743), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n757), .A2(new_n258), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT119), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n993), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT58), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G33), .A2(G41), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT118), .Z(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n406), .C1(G41), .C2(new_n271), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G125), .A2(new_n741), .B1(new_n743), .B2(G137), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n766), .A2(new_n1103), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT120), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1212), .A2(new_n1213), .B1(new_n815), .B2(G132), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n760), .A2(G128), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1211), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n1213), .B2(new_n1212), .C1(new_n994), .C2(new_n765), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT59), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1209), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n751), .A2(G124), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n757), .C2(new_n768), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT121), .Z(new_n1222));
  OAI211_X1 g1022(.A(new_n1207), .B(new_n1210), .C1(new_n1218), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n736), .B1(new_n1223), .B2(new_n737), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1175), .B2(new_n784), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n997), .B2(new_n827), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1198), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1197), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1137), .A2(new_n1231), .A3(new_n956), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n881), .A2(new_n783), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1103), .A2(new_n745), .B1(new_n742), .B2(new_n994), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n271), .B1(new_n750), .B2(new_n1102), .C1(new_n766), .C2(new_n768), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G137), .C2(new_n760), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1205), .B(new_n1236), .C1(new_n406), .C2(new_n765), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n777), .A2(new_n1095), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n742), .A2(new_n519), .B1(new_n745), .B2(new_n450), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n777), .A2(new_n567), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(G283), .C2(new_n760), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n271), .B1(new_n980), .B2(G97), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n987), .A3(new_n1030), .A4(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n750), .A2(new_n478), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1237), .A2(new_n1238), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1245), .A2(new_n737), .B1(new_n259), .B2(new_n828), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1233), .A2(new_n733), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1132), .B2(new_n732), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1232), .A2(new_n1248), .ZN(G381));
  XNOR2_X1  g1049(.A(G375), .B(KEYINPUT124), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1009), .A2(new_n1010), .A3(new_n1074), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1251), .A2(G384), .A3(G381), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1151), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1119), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .A4(new_n1256), .ZN(G407));
  NAND3_X1  g1057(.A1(new_n1250), .A2(new_n665), .A3(new_n1256), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(G213), .A3(new_n1258), .ZN(G409));
  NAND3_X1  g1059(.A1(G378), .A2(new_n1197), .A3(new_n1229), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1189), .A2(new_n956), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1226), .B1(new_n1262), .B2(new_n732), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1255), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(G2897), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1142), .A2(new_n1148), .A3(KEYINPUT60), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1137), .A3(new_n683), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G384), .B(new_n1248), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1231), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1280), .A2(new_n683), .A3(new_n1137), .A4(new_n1274), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1248), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1273), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1248), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1277), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1272), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1271), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1277), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1286), .B2(new_n1277), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1271), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1291), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT126), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1292), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(new_n1007), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1251), .A2(new_n1300), .ZN(new_n1301));
  XOR2_X1   g1101(.A(G393), .B(G396), .Z(new_n1302));
  OR2_X1    g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1074), .A2(new_n975), .A3(new_n1006), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(KEYINPUT127), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1268), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1228), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1264), .B1(new_n1313), .B2(G378), .ZN(new_n1314));
  NOR4_X1   g1114(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1310), .A4(new_n1268), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1299), .B(new_n1307), .C1(new_n1312), .C2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1309), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1321));
  NOR4_X1   g1121(.A1(new_n1314), .A2(KEYINPUT62), .A3(new_n1310), .A4(new_n1268), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1316), .B1(new_n1323), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1256), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1325), .A2(new_n1260), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1290), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1310), .B2(new_n1326), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1307), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1307), .B(new_n1327), .C1(new_n1310), .C2(new_n1326), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(G402));
endmodule


