//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT64), .Z(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n464), .A2(new_n465), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n467), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n466), .B2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n478), .B1(G124), .B2(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n485), .B2(new_n487), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n471), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT4), .B1(new_n467), .B2(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT67), .B1(new_n497), .B2(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT6), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n498), .A2(new_n501), .B1(new_n497), .B2(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(G50), .A3(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT69), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .A3(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n502), .A2(new_n510), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n511), .A2(new_n500), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n505), .A2(new_n514), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n502), .A2(new_n510), .ZN(new_n520));
  AOI211_X1 g095(.A(new_n518), .B(new_n519), .C1(G89), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n498), .A2(new_n501), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n497), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n502), .A2(new_n526), .A3(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND3_X1  g106(.A1(new_n525), .A2(G52), .A3(new_n527), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n507), .A2(new_n509), .A3(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(KEYINPUT72), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G651), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(G90), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n532), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n507), .A2(new_n509), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n520), .A2(G81), .B1(G651), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n525), .A2(G43), .A3(new_n527), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT74), .Z(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n544), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n502), .A2(G91), .A3(new_n510), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n524), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n502), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n563), .A2(new_n564), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n561), .A2(new_n562), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT75), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G299));
  OR2_X1    g148(.A1(new_n505), .A2(new_n514), .ZN(G303));
  OAI21_X1  g149(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  INV_X1    g151(.A(new_n524), .ZN(new_n577));
  AOI22_X1  g152(.A1(G87), .A2(new_n520), .B1(new_n577), .B2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  AOI22_X1  g154(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n500), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n520), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n528), .A2(G47), .ZN(new_n585));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n544), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n520), .A2(G85), .B1(G651), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n512), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n502), .A2(new_n510), .A3(KEYINPUT10), .A4(G92), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n525), .A2(G54), .A3(new_n527), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n500), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  MUX2_X1   g179(.A(G286), .B(G299), .S(new_n604), .Z(G297));
  MUX2_X1   g180(.A(G286), .B(G299), .S(new_n604), .Z(G280));
  INV_X1    g181(.A(G860), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n600), .B1(G559), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT77), .ZN(G148));
  NOR2_X1   g184(.A1(new_n550), .A2(G868), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n600), .A2(G559), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT79), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(G2104), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G2105), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n471), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n467), .A2(G135), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n461), .A2(KEYINPUT80), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT80), .B1(new_n461), .B2(G111), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n624), .A2(G2104), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G123), .B2(new_n482), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n620), .A2(new_n621), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n629), .A2(new_n630), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n622), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(new_n648), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n657), .A2(new_n655), .A3(new_n658), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n655), .A3(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n630), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  AND2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n669), .A2(new_n676), .A3(new_n672), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(G229));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n690));
  NAND2_X1  g265(.A1(G103), .A2(G2104), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G2105), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n467), .A2(G139), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n461), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n699), .B2(G33), .ZN(new_n701));
  INV_X1    g276(.A(G2072), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT91), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n705), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(G1961), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n709));
  INV_X1    g284(.A(G34), .ZN(new_n710));
  AOI21_X1  g285(.A(G29), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G160), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G29), .ZN(new_n715));
  INV_X1    g290(.A(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT94), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT93), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n482), .A2(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT26), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n617), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(new_n699), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n699), .B2(G32), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n718), .B1(G1961), .B2(new_n707), .C1(new_n720), .C2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n701), .A2(new_n702), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n705), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n705), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1966), .ZN(new_n736));
  NAND2_X1  g311(.A1(G164), .A2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G27), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n629), .A2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n742), .B2(KEYINPUT30), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n740), .A2(new_n741), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n729), .A2(new_n720), .ZN(new_n749));
  INV_X1    g324(.A(new_n715), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n750), .A2(G2084), .B1(new_n739), .B2(new_n738), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n733), .A2(new_n736), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n708), .A2(new_n731), .A3(new_n732), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n705), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n699), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n699), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT29), .Z(new_n763));
  OAI21_X1  g338(.A(new_n759), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n760), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n705), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n550), .B2(new_n705), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1341), .Z(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT89), .Z(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n600), .B2(new_n705), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n699), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(G116), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n616), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n467), .A2(G140), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G128), .B2(new_n482), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n699), .ZN(new_n783));
  INV_X1    g358(.A(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n767), .A2(new_n770), .A3(new_n774), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n765), .B2(KEYINPUT97), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n755), .A2(new_n766), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n705), .A2(G6), .ZN(new_n789));
  INV_X1    g364(.A(G305), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n705), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1981), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G1981), .ZN(new_n794));
  NOR2_X1   g369(.A1(G166), .A2(new_n705), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n705), .B2(G22), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n705), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(G288), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n705), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT33), .B(G1976), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n797), .A2(G1971), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  INV_X1    g379(.A(new_n800), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n796), .A2(new_n804), .B1(new_n805), .B2(new_n801), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n793), .A2(new_n794), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n699), .A2(G25), .ZN(new_n810));
  NOR2_X1   g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT86), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT87), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n482), .A2(G119), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n467), .A2(G131), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT88), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n810), .B1(new_n818), .B2(new_n699), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n705), .A2(G24), .ZN(new_n824));
  INV_X1    g399(.A(G290), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n825), .B2(new_n705), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1986), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n808), .A2(new_n809), .A3(new_n822), .A4(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT36), .Z(new_n830));
  NOR2_X1   g405(.A1(new_n788), .A2(new_n830), .ZN(G311));
  OR2_X1    g406(.A1(new_n788), .A2(new_n830), .ZN(G150));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n544), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n520), .A2(G93), .B1(G651), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n525), .A2(G55), .A3(new_n527), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n601), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n549), .A2(new_n838), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n547), .A2(new_n836), .A3(new_n548), .A4(new_n837), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n843), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n607), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n840), .B1(new_n849), .B2(new_n850), .ZN(G145));
  OR2_X1    g426(.A1(new_n817), .A2(new_n619), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n817), .A2(new_n619), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n467), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n858), .B1(G130), .B2(new_n482), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n852), .A2(new_n859), .A3(new_n853), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(KEYINPUT100), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n494), .A2(new_n495), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n726), .B(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n782), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n782), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n697), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n696), .A3(new_n868), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n869), .B2(new_n870), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n864), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n869), .A2(new_n870), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n876), .A2(new_n863), .A3(new_n871), .A4(new_n873), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n714), .B(G162), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n629), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT101), .Z(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT102), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n876), .A2(new_n871), .A3(new_n873), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n861), .A2(new_n862), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n879), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g468(.A1(new_n838), .A2(new_n604), .ZN(new_n894));
  XNOR2_X1  g469(.A(G290), .B(new_n790), .ZN(new_n895));
  XNOR2_X1  g470(.A(G166), .B(G288), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  XOR2_X1   g473(.A(new_n611), .B(new_n846), .Z(new_n899));
  NAND3_X1  g474(.A1(new_n600), .A2(new_n569), .A3(new_n572), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n600), .B1(new_n572), .B2(new_n569), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT41), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(G299), .A2(new_n601), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n600), .A2(new_n569), .A3(new_n572), .A4(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n899), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n901), .A2(new_n902), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n899), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n898), .B1(KEYINPUT104), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(KEYINPUT104), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n898), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n894), .B1(new_n915), .B2(new_n604), .ZN(G331));
  XNOR2_X1  g491(.A(G331), .B(KEYINPUT105), .ZN(G295));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g493(.A1(G301), .A2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n532), .A2(new_n539), .A3(new_n540), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n844), .A3(new_n845), .ZN(new_n923));
  AND4_X1   g498(.A1(new_n548), .A2(new_n547), .A3(new_n836), .A4(new_n837), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n548), .A2(new_n547), .B1(new_n836), .B2(new_n837), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n919), .B(new_n921), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G286), .ZN(new_n928));
  INV_X1    g503(.A(new_n911), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n926), .A3(G168), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n897), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n909), .A2(new_n903), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n930), .B2(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  AOI21_X1  g511(.A(G168), .B1(new_n923), .B2(new_n926), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n903), .B(new_n909), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n931), .A4(new_n897), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n905), .B1(new_n928), .B2(new_n930), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n897), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n911), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n941), .A2(new_n942), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n897), .B1(new_n938), .B2(new_n931), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(G37), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n942), .B1(new_n941), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n952), .B2(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n954), .B(new_n942), .C1(new_n941), .C2(new_n951), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n918), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n941), .A2(new_n948), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n918), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n941), .A2(new_n942), .A3(new_n951), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n956), .B(new_n965), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n865), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT112), .B(G40), .Z(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n782), .B(G2067), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n727), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1996), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n974), .A2(KEYINPUT46), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT46), .B1(new_n974), .B2(new_n978), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT47), .Z(new_n982));
  NOR2_X1   g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT113), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(new_n974), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT48), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n727), .A2(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n726), .A2(G1996), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n976), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n974), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n817), .A2(new_n820), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n817), .A2(new_n820), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n974), .A3(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n985), .A2(KEYINPUT48), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n986), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n990), .A2(new_n818), .A3(new_n820), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n782), .A2(new_n784), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n974), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n982), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT49), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n969), .ZN(new_n1004));
  AND2_X1   g579(.A1(G160), .A2(new_n972), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n1002), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1007), .B1(G1976), .B2(new_n799), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(KEYINPUT115), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT115), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1010), .B(new_n1013), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n973), .B1(new_n1004), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n971), .B(new_n1005), .C1(new_n1027), .C2(new_n969), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1026), .A2(G2090), .B1(new_n1029), .B2(G1971), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT55), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1019), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1010), .A2(new_n1014), .A3(new_n799), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT116), .A3(new_n1001), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n1036), .B2(new_n1001), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1007), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n760), .B1(new_n804), .B2(new_n1028), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1033), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1034), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1019), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1018), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1016), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT117), .A3(new_n1010), .A4(new_n1013), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1045), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n973), .B1(new_n1027), .B2(new_n969), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n969), .B2(new_n970), .ZN(new_n1053));
  INV_X1    g628(.A(G1966), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n716), .B(new_n1021), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1043), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1057), .A2(G168), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT63), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1034), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1019), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1040), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT53), .B1(new_n1029), .B2(new_n739), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(KEYINPUT126), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT126), .ZN(new_n1067));
  INV_X1    g642(.A(G1961), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1026), .A2(KEYINPUT121), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1070), .B(new_n1021), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n739), .A2(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1053), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G168), .A2(new_n1043), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n1057), .A2(KEYINPUT125), .A3(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1076), .B(KEYINPUT124), .Z(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT51), .B1(new_n1079), .B2(new_n1057), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT125), .B1(new_n1057), .B2(new_n1077), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1076), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(KEYINPUT62), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT62), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1086));
  OAI211_X1 g661(.A(G171), .B(new_n1075), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n570), .A2(KEYINPUT57), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(new_n563), .C1(KEYINPUT119), .C2(KEYINPUT57), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n563), .A2(KEYINPUT119), .B1(new_n570), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT118), .B1(new_n567), .B2(new_n568), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1093), .B2(KEYINPUT57), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT120), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT56), .B(G2072), .Z(new_n1096));
  OAI22_X1  g671(.A1(new_n1041), .A2(G1956), .B1(new_n1028), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1006), .A2(G2067), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1072), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(new_n600), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1006), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT122), .B(G1996), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1028), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n550), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(KEYINPUT123), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1110), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n600), .B1(new_n1101), .B2(KEYINPUT60), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1095), .B(new_n1097), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1104), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G301), .B(KEYINPUT54), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n971), .B1(new_n1027), .B2(new_n969), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G40), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n714), .A2(new_n1124), .A3(new_n1074), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1075), .A2(new_n1121), .B1(new_n1073), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1087), .B1(new_n1120), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1064), .B1(new_n1130), .B2(new_n1051), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n984), .B1(G1986), .B2(G290), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n994), .B1(new_n1132), .B2(new_n975), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1000), .B1(new_n1131), .B2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g709(.A1(G227), .A2(new_n459), .ZN(new_n1136));
  NAND4_X1  g710(.A1(new_n687), .A2(new_n653), .A3(new_n688), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g711(.A(new_n1137), .B1(new_n885), .B2(new_n891), .ZN(new_n1138));
  OAI211_X1 g712(.A(new_n1138), .B(KEYINPUT127), .C1(new_n955), .C2(new_n953), .ZN(new_n1139));
  INV_X1    g713(.A(new_n1139), .ZN(new_n1140));
  OR2_X1    g714(.A1(new_n953), .A2(new_n955), .ZN(new_n1141));
  AOI21_X1  g715(.A(KEYINPUT127), .B1(new_n1141), .B2(new_n1138), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1142), .ZN(G308));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1138), .ZN(G225));
endmodule


