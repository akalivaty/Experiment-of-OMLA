

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744;

  NAND2_X1 U367 ( .A1(n346), .A2(n345), .ZN(n521) );
  INV_X1 U368 ( .A(n664), .ZN(n345) );
  INV_X1 U369 ( .A(n651), .ZN(n346) );
  AND2_X2 U370 ( .A1(n385), .A2(n386), .ZN(n384) );
  INV_X1 U371 ( .A(G953), .ZN(n734) );
  NOR2_X1 U372 ( .A1(n511), .A2(n503), .ZN(n504) );
  XNOR2_X2 U373 ( .A(n549), .B(n548), .ZN(n594) );
  AND2_X2 U374 ( .A1(n565), .A2(n672), .ZN(n548) );
  XNOR2_X2 U375 ( .A(n365), .B(n531), .ZN(n721) );
  NAND2_X2 U376 ( .A1(n370), .A2(n369), .ZN(n365) );
  XNOR2_X2 U377 ( .A(n493), .B(n492), .ZN(n551) );
  XNOR2_X2 U378 ( .A(n514), .B(KEYINPUT31), .ZN(n664) );
  XNOR2_X2 U379 ( .A(n469), .B(G472), .ZN(n512) );
  XNOR2_X1 U380 ( .A(G143), .B(G128), .ZN(n441) );
  XNOR2_X1 U381 ( .A(G101), .B(KEYINPUT72), .ZN(n397) );
  AND2_X1 U382 ( .A1(n372), .A2(n530), .ZN(n371) );
  AND2_X1 U383 ( .A1(n544), .A2(n543), .ZN(n565) );
  AND2_X1 U384 ( .A1(n494), .A2(n503), .ZN(n393) );
  XNOR2_X1 U385 ( .A(n606), .B(n605), .ZN(n607) );
  XOR2_X1 U386 ( .A(KEYINPUT122), .B(n633), .Z(n634) );
  XNOR2_X1 U387 ( .A(n441), .B(G134), .ZN(n455) );
  XNOR2_X1 U388 ( .A(n397), .B(n399), .ZN(n381) );
  XNOR2_X1 U389 ( .A(G119), .B(G113), .ZN(n398) );
  XNOR2_X1 U390 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X2 U391 ( .A(n428), .B(KEYINPUT10), .ZN(n731) );
  OR2_X2 U392 ( .A1(n604), .A2(G902), .ZN(n357) );
  NOR2_X1 U393 ( .A1(n670), .A2(n505), .ZN(n506) );
  XNOR2_X1 U394 ( .A(n499), .B(n368), .ZN(n374) );
  INV_X1 U395 ( .A(KEYINPUT64), .ZN(n368) );
  NAND2_X1 U396 ( .A1(n392), .A2(n347), .ZN(n383) );
  XNOR2_X1 U397 ( .A(n459), .B(n458), .ZN(n732) );
  XNOR2_X1 U398 ( .A(n455), .B(G137), .ZN(n459) );
  XOR2_X1 U399 ( .A(G146), .B(G125), .Z(n427) );
  XOR2_X1 U400 ( .A(G140), .B(KEYINPUT79), .Z(n472) );
  XNOR2_X1 U401 ( .A(n717), .B(KEYINPUT73), .ZN(n476) );
  XNOR2_X1 U402 ( .A(n502), .B(KEYINPUT74), .ZN(n511) );
  INV_X1 U403 ( .A(n553), .ZN(n539) );
  XNOR2_X1 U404 ( .A(n357), .B(n356), .ZN(n686) );
  XNOR2_X1 U405 ( .A(G469), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U406 ( .A(n732), .B(G146), .ZN(n379) );
  NAND2_X1 U407 ( .A1(n424), .A2(n396), .ZN(n426) );
  NOR2_X1 U408 ( .A1(n511), .A2(n541), .ZN(n694) );
  NAND2_X1 U409 ( .A1(KEYINPUT84), .A2(n390), .ZN(n389) );
  INV_X1 U410 ( .A(KEYINPUT44), .ZN(n390) );
  INV_X1 U411 ( .A(G237), .ZN(n411) );
  AND2_X1 U412 ( .A1(n582), .A2(n581), .ZN(n585) );
  NOR2_X1 U413 ( .A1(n374), .A2(n373), .ZN(n376) );
  XNOR2_X1 U414 ( .A(KEYINPUT70), .B(G131), .ZN(n457) );
  XOR2_X1 U415 ( .A(G122), .B(G104), .Z(n430) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT89), .ZN(n405) );
  XOR2_X1 U417 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n456) );
  XOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT18), .Z(n402) );
  INV_X1 U419 ( .A(n357), .ZN(n478) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n462) );
  XOR2_X1 U421 ( .A(G116), .B(KEYINPUT5), .Z(n461) );
  XNOR2_X1 U422 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U423 ( .A(G101), .B(G107), .ZN(n473) );
  NOR2_X1 U424 ( .A1(n587), .A2(n541), .ZN(n542) );
  INV_X1 U425 ( .A(KEYINPUT92), .ZN(n358) );
  BUF_X1 U426 ( .A(n512), .Z(n692) );
  AND2_X2 U427 ( .A1(n382), .A2(n603), .ZN(n712) );
  XNOR2_X1 U428 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U429 ( .A(n610), .B(KEYINPUT86), .ZN(n643) );
  AND2_X1 U430 ( .A1(n495), .A2(n503), .ZN(n523) );
  NOR2_X1 U431 ( .A1(n624), .A2(n716), .ZN(n625) );
  XNOR2_X1 U432 ( .A(n395), .B(n623), .ZN(n624) );
  XNOR2_X1 U433 ( .A(n711), .B(n366), .ZN(G75) );
  XNOR2_X1 U434 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n366) );
  AND2_X1 U435 ( .A1(n525), .A2(KEYINPUT84), .ZN(n347) );
  XOR2_X1 U436 ( .A(G104), .B(KEYINPUT76), .Z(n348) );
  OR2_X1 U437 ( .A1(n692), .A2(n532), .ZN(n349) );
  AND2_X1 U438 ( .A1(n557), .A2(n682), .ZN(n350) );
  XOR2_X1 U439 ( .A(KEYINPUT47), .B(n564), .Z(n351) );
  INV_X1 U440 ( .A(n686), .ZN(n500) );
  XOR2_X1 U441 ( .A(n417), .B(KEYINPUT19), .Z(n352) );
  XNOR2_X1 U442 ( .A(n379), .B(n477), .ZN(n604) );
  INV_X1 U443 ( .A(KEYINPUT84), .ZN(n526) );
  INV_X1 U444 ( .A(KEYINPUT83), .ZN(n373) );
  AND2_X1 U445 ( .A1(n603), .A2(G210), .ZN(n353) );
  AND2_X1 U446 ( .A1(n526), .A2(KEYINPUT44), .ZN(n354) );
  NAND2_X1 U447 ( .A1(n598), .A2(KEYINPUT2), .ZN(n355) );
  NOR2_X2 U448 ( .A1(n349), .A2(n505), .ZN(n651) );
  XNOR2_X2 U449 ( .A(n513), .B(n358), .ZN(n505) );
  OR2_X2 U450 ( .A1(n359), .A2(n476), .ZN(n363) );
  XNOR2_X1 U451 ( .A(n348), .B(G110), .ZN(n717) );
  XNOR2_X1 U452 ( .A(n466), .B(n380), .ZN(n359) );
  XNOR2_X2 U453 ( .A(n442), .B(KEYINPUT16), .ZN(n380) );
  XNOR2_X2 U454 ( .A(n381), .B(n398), .ZN(n466) );
  OR2_X1 U455 ( .A1(n377), .A2(KEYINPUT83), .ZN(n369) );
  XNOR2_X1 U456 ( .A(n478), .B(G469), .ZN(n360) );
  XNOR2_X1 U457 ( .A(n466), .B(n380), .ZN(n361) );
  NAND2_X1 U458 ( .A1(n361), .A2(n476), .ZN(n362) );
  NAND2_X1 U459 ( .A1(n362), .A2(n363), .ZN(n410) );
  NOR2_X2 U460 ( .A1(n551), .A2(n501), .ZN(n685) );
  XNOR2_X1 U461 ( .A(G143), .B(G128), .ZN(n364) );
  NAND2_X1 U462 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U463 ( .A1(n377), .A2(n376), .ZN(n375) );
  XNOR2_X2 U464 ( .A(n367), .B(n454), .ZN(n495) );
  NAND2_X1 U465 ( .A1(n350), .A2(n513), .ZN(n367) );
  XNOR2_X2 U466 ( .A(n426), .B(n425), .ZN(n513) );
  AND2_X2 U467 ( .A1(n375), .A2(n371), .ZN(n370) );
  NAND2_X1 U468 ( .A1(n384), .A2(n383), .ZN(n377) );
  NAND2_X2 U469 ( .A1(n545), .A2(n671), .ZN(n575) );
  XNOR2_X1 U470 ( .A(n379), .B(n467), .ZN(n628) );
  XNOR2_X2 U471 ( .A(n400), .B(G107), .ZN(n442) );
  INV_X1 U472 ( .A(n424), .ZN(n561) );
  XNOR2_X2 U473 ( .A(n575), .B(n352), .ZN(n424) );
  XNOR2_X2 U474 ( .A(n413), .B(n412), .ZN(n545) );
  NAND2_X1 U475 ( .A1(n527), .A2(n354), .ZN(n385) );
  AND2_X2 U476 ( .A1(n524), .A2(n616), .ZN(n525) );
  AND2_X1 U477 ( .A1(n382), .A2(n669), .ZN(n709) );
  NAND2_X1 U478 ( .A1(n382), .A2(n353), .ZN(n395) );
  XNOR2_X2 U479 ( .A(n599), .B(n355), .ZN(n382) );
  NAND2_X1 U480 ( .A1(n387), .A2(n388), .ZN(n386) );
  NAND2_X1 U481 ( .A1(n391), .A2(KEYINPUT84), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n525), .A2(n389), .ZN(n388) );
  INV_X1 U483 ( .A(n525), .ZN(n391) );
  INV_X1 U484 ( .A(n527), .ZN(n392) );
  XNOR2_X2 U485 ( .A(n510), .B(KEYINPUT35), .ZN(n527) );
  NAND2_X1 U486 ( .A1(n495), .A2(n393), .ZN(n394) );
  NAND2_X1 U487 ( .A1(n618), .A2(n614), .ZN(n528) );
  XNOR2_X2 U488 ( .A(n394), .B(KEYINPUT32), .ZN(n618) );
  AND2_X1 U489 ( .A1(n701), .A2(n423), .ZN(n396) );
  INV_X1 U490 ( .A(n667), .ZN(n579) );
  XNOR2_X1 U491 ( .A(n427), .B(n402), .ZN(n403) );
  NOR2_X1 U492 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U493 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U494 ( .A(n476), .B(n475), .ZN(n477) );
  AND2_X1 U495 ( .A1(n540), .A2(n539), .ZN(n544) );
  BUF_X1 U496 ( .A(n361), .Z(n718) );
  XNOR2_X2 U497 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X2 U498 ( .A(G122), .B(G116), .ZN(n400) );
  NAND2_X1 U499 ( .A1(G224), .A2(n734), .ZN(n401) );
  XNOR2_X1 U500 ( .A(n401), .B(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U501 ( .A(n364), .B(n405), .ZN(n406) );
  XNOR2_X1 U502 ( .A(n456), .B(n406), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U504 ( .A(n410), .B(n409), .ZN(n619) );
  XNOR2_X1 U505 ( .A(KEYINPUT15), .B(G902), .ZN(n601) );
  NAND2_X1 U506 ( .A1(n619), .A2(n601), .ZN(n413) );
  INV_X1 U507 ( .A(G902), .ZN(n468) );
  NAND2_X1 U508 ( .A1(n468), .A2(n411), .ZN(n414) );
  AND2_X1 U509 ( .A1(n414), .A2(G210), .ZN(n412) );
  NAND2_X1 U510 ( .A1(n414), .A2(G214), .ZN(n416) );
  INV_X1 U511 ( .A(KEYINPUT91), .ZN(n415) );
  XNOR2_X1 U512 ( .A(n416), .B(n415), .ZN(n671) );
  INV_X1 U513 ( .A(KEYINPUT66), .ZN(n417) );
  NAND2_X1 U514 ( .A1(G237), .A2(G234), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n418), .B(KEYINPUT14), .ZN(n701) );
  AND2_X1 U516 ( .A1(n734), .A2(G952), .ZN(n536) );
  INV_X1 U517 ( .A(n536), .ZN(n422) );
  INV_X1 U518 ( .A(G898), .ZN(n420) );
  NAND2_X1 U519 ( .A1(G953), .A2(G902), .ZN(n533) );
  INV_X1 U520 ( .A(n533), .ZN(n419) );
  NAND2_X1 U521 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND2_X1 U522 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U523 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n425) );
  XNOR2_X1 U524 ( .A(G140), .B(n427), .ZN(n428) );
  XNOR2_X1 U525 ( .A(G143), .B(G113), .ZN(n429) );
  XNOR2_X1 U526 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U527 ( .A(n731), .B(n431), .ZN(n438) );
  XOR2_X1 U528 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n433) );
  NAND2_X1 U529 ( .A1(G214), .A2(n462), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U531 ( .A(KEYINPUT11), .B(n434), .ZN(n436) );
  INV_X1 U532 ( .A(n457), .ZN(n435) );
  XOR2_X1 U533 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U534 ( .A(n438), .B(n437), .ZN(n640) );
  NOR2_X1 U535 ( .A1(G902), .A2(n640), .ZN(n440) );
  XNOR2_X1 U536 ( .A(KEYINPUT13), .B(G475), .ZN(n439) );
  XNOR2_X1 U537 ( .A(n440), .B(n439), .ZN(n519) );
  XOR2_X1 U538 ( .A(n455), .B(n442), .Z(n448) );
  XOR2_X1 U539 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n446) );
  NAND2_X1 U540 ( .A1(n734), .A2(G234), .ZN(n444) );
  XNOR2_X1 U541 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n443) );
  XNOR2_X1 U542 ( .A(n444), .B(n443), .ZN(n484) );
  NAND2_X1 U543 ( .A1(G217), .A2(n484), .ZN(n445) );
  XNOR2_X1 U544 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U545 ( .A(n448), .B(n447), .ZN(n633) );
  NOR2_X1 U546 ( .A1(G902), .A2(n633), .ZN(n449) );
  XOR2_X1 U547 ( .A(G478), .B(n449), .Z(n516) );
  NOR2_X1 U548 ( .A1(n519), .A2(n516), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n450), .B(KEYINPUT98), .ZN(n557) );
  NAND2_X1 U550 ( .A1(G234), .A2(n601), .ZN(n451) );
  XNOR2_X1 U551 ( .A(KEYINPUT20), .B(n451), .ZN(n489) );
  AND2_X1 U552 ( .A1(n489), .A2(G221), .ZN(n453) );
  INV_X1 U553 ( .A(KEYINPUT21), .ZN(n452) );
  XNOR2_X1 U554 ( .A(n453), .B(n452), .ZN(n501) );
  INV_X1 U555 ( .A(n501), .ZN(n682) );
  INV_X1 U556 ( .A(KEYINPUT22), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT75), .ZN(n460) );
  XNOR2_X1 U559 ( .A(n461), .B(n460), .ZN(n464) );
  NAND2_X1 U560 ( .A1(n462), .A2(G210), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U562 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U563 ( .A1(n628), .A2(n468), .ZN(n469) );
  INV_X1 U564 ( .A(KEYINPUT6), .ZN(n470) );
  XNOR2_X1 U565 ( .A(n512), .B(n470), .ZN(n569) );
  INV_X1 U566 ( .A(n569), .ZN(n503) );
  NAND2_X1 U567 ( .A1(G227), .A2(n734), .ZN(n471) );
  XNOR2_X1 U568 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U569 ( .A(n500), .B(KEYINPUT85), .ZN(n577) );
  XOR2_X1 U570 ( .A(G110), .B(G119), .Z(n480) );
  XNOR2_X1 U571 ( .A(G128), .B(G137), .ZN(n479) );
  XNOR2_X1 U572 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U573 ( .A(n731), .B(n481), .ZN(n488) );
  XNOR2_X1 U574 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n482) );
  XNOR2_X1 U575 ( .A(n482), .B(KEYINPUT93), .ZN(n483) );
  XOR2_X1 U576 ( .A(KEYINPUT94), .B(n483), .Z(n486) );
  NAND2_X1 U577 ( .A1(G221), .A2(n484), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n488), .B(n487), .ZN(n713) );
  NOR2_X1 U580 ( .A1(n713), .A2(G902), .ZN(n493) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT25), .Z(n491) );
  NAND2_X1 U582 ( .A1(n489), .A2(G217), .ZN(n490) );
  XNOR2_X1 U583 ( .A(n491), .B(n490), .ZN(n492) );
  AND2_X1 U584 ( .A1(n577), .A2(n551), .ZN(n494) );
  INV_X1 U585 ( .A(n495), .ZN(n498) );
  INV_X1 U586 ( .A(n551), .ZN(n683) );
  NOR2_X1 U587 ( .A1(n692), .A2(n683), .ZN(n496) );
  NAND2_X1 U588 ( .A1(n496), .A2(n500), .ZN(n497) );
  OR2_X1 U589 ( .A1(n498), .A2(n497), .ZN(n614) );
  NAND2_X1 U590 ( .A1(n528), .A2(KEYINPUT44), .ZN(n499) );
  NAND2_X1 U591 ( .A1(n686), .A2(n685), .ZN(n502) );
  XNOR2_X1 U592 ( .A(n504), .B(KEYINPUT33), .ZN(n670) );
  XNOR2_X1 U593 ( .A(n506), .B(KEYINPUT34), .ZN(n509) );
  NAND2_X1 U594 ( .A1(n516), .A2(n519), .ZN(n567) );
  INV_X1 U595 ( .A(KEYINPUT80), .ZN(n507) );
  XNOR2_X1 U596 ( .A(n567), .B(n507), .ZN(n508) );
  NAND2_X1 U597 ( .A1(n509), .A2(n508), .ZN(n510) );
  INV_X1 U598 ( .A(n512), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n694), .A2(n513), .ZN(n514) );
  INV_X1 U600 ( .A(n685), .ZN(n515) );
  OR2_X1 U601 ( .A1(n360), .A2(n515), .ZN(n532) );
  INV_X1 U602 ( .A(n516), .ZN(n518) );
  NOR2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n517) );
  XOR2_X1 U604 ( .A(KEYINPUT97), .B(n517), .Z(n663) );
  NAND2_X1 U605 ( .A1(n519), .A2(n518), .ZN(n572) );
  INV_X1 U606 ( .A(n572), .ZN(n520) );
  NOR2_X1 U607 ( .A1(n663), .A2(n520), .ZN(n677) );
  INV_X1 U608 ( .A(n677), .ZN(n563) );
  NAND2_X1 U609 ( .A1(n521), .A2(n563), .ZN(n524) );
  AND2_X1 U610 ( .A1(n500), .A2(n683), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n616) );
  NOR2_X1 U612 ( .A1(n528), .A2(KEYINPUT44), .ZN(n529) );
  NAND2_X1 U613 ( .A1(n392), .A2(n529), .ZN(n530) );
  INV_X1 U614 ( .A(KEYINPUT45), .ZN(n531) );
  XNOR2_X1 U615 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n549) );
  INV_X1 U616 ( .A(n532), .ZN(n540) );
  NOR2_X1 U617 ( .A1(G900), .A2(n533), .ZN(n534) );
  NAND2_X1 U618 ( .A1(n701), .A2(n534), .ZN(n535) );
  XOR2_X1 U619 ( .A(KEYINPUT100), .B(n535), .Z(n538) );
  AND2_X1 U620 ( .A1(n536), .A2(n701), .ZN(n537) );
  NOR2_X1 U621 ( .A1(n538), .A2(n537), .ZN(n553) );
  INV_X1 U622 ( .A(n671), .ZN(n587) );
  XNOR2_X1 U623 ( .A(KEYINPUT30), .B(n542), .ZN(n543) );
  BUF_X1 U624 ( .A(n545), .Z(n546) );
  INV_X1 U625 ( .A(KEYINPUT38), .ZN(n547) );
  XNOR2_X1 U626 ( .A(n546), .B(n547), .ZN(n672) );
  NOR2_X1 U627 ( .A1(n572), .A2(n594), .ZN(n550) );
  XNOR2_X1 U628 ( .A(n550), .B(KEYINPUT40), .ZN(n742) );
  NAND2_X1 U629 ( .A1(n551), .A2(n682), .ZN(n552) );
  NOR2_X1 U630 ( .A1(n553), .A2(n552), .ZN(n570) );
  AND2_X1 U631 ( .A1(n692), .A2(n570), .ZN(n554) );
  XNOR2_X1 U632 ( .A(KEYINPUT28), .B(n554), .ZN(n556) );
  INV_X1 U633 ( .A(n360), .ZN(n555) );
  NAND2_X1 U634 ( .A1(n556), .A2(n555), .ZN(n562) );
  NAND2_X1 U635 ( .A1(n672), .A2(n671), .ZN(n676) );
  INV_X1 U636 ( .A(n557), .ZN(n675) );
  NOR2_X1 U637 ( .A1(n676), .A2(n675), .ZN(n558) );
  XNOR2_X1 U638 ( .A(n558), .B(KEYINPUT41), .ZN(n704) );
  NOR2_X1 U639 ( .A1(n562), .A2(n704), .ZN(n559) );
  XNOR2_X1 U640 ( .A(n559), .B(KEYINPUT42), .ZN(n743) );
  NOR2_X2 U641 ( .A1(n742), .A2(n743), .ZN(n560) );
  XNOR2_X1 U642 ( .A(n560), .B(KEYINPUT46), .ZN(n582) );
  NOR2_X1 U643 ( .A1(n562), .A2(n561), .ZN(n658) );
  NAND2_X1 U644 ( .A1(n658), .A2(n563), .ZN(n564) );
  INV_X1 U645 ( .A(n565), .ZN(n566) );
  NOR2_X1 U646 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U647 ( .A1(n568), .A2(n546), .ZN(n613) );
  NAND2_X1 U648 ( .A1(n351), .A2(n613), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U650 ( .A(KEYINPUT101), .B(n571), .ZN(n573) );
  XNOR2_X1 U651 ( .A(KEYINPUT99), .B(n572), .ZN(n661) );
  NAND2_X1 U652 ( .A1(n573), .A2(n661), .ZN(n574) );
  XNOR2_X1 U653 ( .A(KEYINPUT102), .B(n574), .ZN(n586) );
  NOR2_X1 U654 ( .A1(n586), .A2(n575), .ZN(n576) );
  XNOR2_X1 U655 ( .A(n576), .B(KEYINPUT36), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n667) );
  INV_X1 U657 ( .A(KEYINPUT71), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT48), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n585), .B(n584), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n500), .A2(n588), .ZN(n589) );
  XNOR2_X1 U662 ( .A(KEYINPUT103), .B(n589), .ZN(n590) );
  XOR2_X1 U663 ( .A(n590), .B(KEYINPUT43), .Z(n592) );
  INV_X1 U664 ( .A(n546), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n617) );
  INV_X1 U666 ( .A(n663), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n668) );
  INV_X1 U668 ( .A(n668), .ZN(n595) );
  AND2_X1 U669 ( .A1(n617), .A2(n595), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n730) );
  NOR2_X2 U671 ( .A1(n721), .A2(n730), .ZN(n599) );
  INV_X1 U672 ( .A(KEYINPUT77), .ZN(n598) );
  INV_X1 U673 ( .A(KEYINPUT2), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n600), .A2(KEYINPUT77), .ZN(n669) );
  INV_X1 U675 ( .A(n601), .ZN(n602) );
  AND2_X1 U676 ( .A1(n669), .A2(n602), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n712), .A2(G469), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT57), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n608), .B(n607), .ZN(n611) );
  INV_X1 U681 ( .A(G952), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n609), .A2(G953), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n643), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT119), .ZN(G54) );
  XNOR2_X1 U685 ( .A(n613), .B(G143), .ZN(G45) );
  XNOR2_X1 U686 ( .A(n614), .B(G110), .ZN(G12) );
  XNOR2_X1 U687 ( .A(G101), .B(KEYINPUT106), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G3) );
  XNOR2_X1 U689 ( .A(n617), .B(G140), .ZN(G42) );
  XOR2_X1 U690 ( .A(G122), .B(n527), .Z(G24) );
  XNOR2_X1 U691 ( .A(n618), .B(G119), .ZN(G21) );
  BUF_X1 U692 ( .A(n619), .Z(n620) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(KEYINPUT54), .Z(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT55), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n620), .B(n622), .ZN(n623) );
  INV_X1 U696 ( .A(n643), .ZN(n716) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U698 ( .A1(n712), .A2(G472), .ZN(n630) );
  XOR2_X1 U699 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(KEYINPUT62), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n631), .A2(n643), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U704 ( .A1(n712), .A2(G478), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n636), .A2(n643), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U708 ( .A1(n712), .A2(G475), .ZN(n642) );
  XOR2_X1 U709 ( .A(KEYINPUT65), .B(KEYINPUT120), .Z(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT59), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U713 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(G60) );
  XOR2_X1 U715 ( .A(G104), .B(KEYINPUT107), .Z(n648) );
  NAND2_X1 U716 ( .A1(n651), .A2(n661), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n648), .B(n647), .ZN(G6) );
  XOR2_X1 U718 ( .A(KEYINPUT110), .B(KEYINPUT27), .Z(n650) );
  XNOR2_X1 U719 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n650), .B(n649), .ZN(n655) );
  XOR2_X1 U721 ( .A(G107), .B(KEYINPUT26), .Z(n653) );
  NAND2_X1 U722 ( .A1(n651), .A2(n663), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G9) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .Z(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n663), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(G30) );
  XOR2_X1 U728 ( .A(G146), .B(KEYINPUT111), .Z(n660) );
  NAND2_X1 U729 ( .A1(n658), .A2(n661), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n664), .A2(n661), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(G113), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n665), .B(G116), .ZN(G18) );
  XOR2_X1 U735 ( .A(G125), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(G27) );
  XOR2_X1 U737 ( .A(G134), .B(n668), .Z(G36) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT114), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT115), .B(n680), .Z(n681) );
  NOR2_X1 U744 ( .A1(n670), .A2(n681), .ZN(n699) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U746 ( .A(KEYINPUT49), .B(n684), .ZN(n690) );
  OR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U748 ( .A(n687), .B(KEYINPUT112), .ZN(n688) );
  XNOR2_X1 U749 ( .A(KEYINPUT50), .B(n688), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n695), .B(KEYINPUT51), .ZN(n696) );
  XNOR2_X1 U754 ( .A(KEYINPUT113), .B(n696), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n704), .A2(n697), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U757 ( .A(KEYINPUT52), .B(n700), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n701), .A2(G952), .ZN(n702) );
  OR2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n670), .A2(n704), .ZN(n705) );
  XOR2_X1 U761 ( .A(KEYINPUT116), .B(n705), .Z(n706) );
  NAND2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U764 ( .A1(n734), .A2(n710), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n712), .A2(G217), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(G66) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U769 ( .A1(G898), .A2(n734), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n729) );
  BUF_X1 U771 ( .A(n721), .Z(n722) );
  NOR2_X1 U772 ( .A1(n722), .A2(G953), .ZN(n723) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(n723), .Z(n727) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n724) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U776 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U777 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(G69) );
  XNOR2_X1 U779 ( .A(KEYINPUT125), .B(n730), .ZN(n733) );
  XOR2_X1 U780 ( .A(n732), .B(n731), .Z(n737) );
  XOR2_X1 U781 ( .A(n733), .B(n737), .Z(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U783 ( .A(n736), .B(KEYINPUT126), .ZN(n741) );
  XNOR2_X1 U784 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n741), .A2(n740), .ZN(G72) );
  XOR2_X1 U788 ( .A(n742), .B(G131), .Z(G33) );
  XNOR2_X1 U789 ( .A(G137), .B(KEYINPUT127), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(G39) );
endmodule

