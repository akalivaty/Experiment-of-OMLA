//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n203), .C2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NOR2_X1   g0032(.A1(G58), .A2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n228), .B1(new_n232), .B2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  INV_X1    g0043(.A(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n229), .ZN(new_n257));
  INV_X1    g0057(.A(G20), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n260), .A2(new_n213), .B1(new_n258), .B2(G68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n215), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n257), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(new_n264), .B(KEYINPUT11), .Z(new_n265));
  INV_X1    g0065(.A(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G1), .B2(new_n258), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n208), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n258), .A3(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n208), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT12), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n265), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(G1), .B(G13), .C1(new_n259), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G238), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n214), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n219), .A2(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n282), .B(new_n285), .C1(new_n278), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n289), .A3(new_n290), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n278), .B1(new_n296), .B2(new_n286), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n282), .A4(new_n285), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n276), .B1(new_n301), .B2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI211_X1 g0103(.A(KEYINPUT14), .B(new_n303), .C1(new_n295), .C2(new_n300), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n295), .A2(G179), .A3(new_n300), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT70), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n297), .A2(new_n284), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n299), .B1(new_n308), .B2(new_n282), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n278), .A2(new_n280), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n209), .ZN(new_n311));
  NOR4_X1   g0111(.A1(new_n297), .A2(new_n311), .A3(KEYINPUT13), .A4(new_n284), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n301), .A2(new_n276), .A3(G169), .ZN(new_n315));
  AND4_X1   g0115(.A1(KEYINPUT70), .A2(new_n314), .A3(new_n306), .A4(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n275), .B1(new_n307), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n288), .A2(G222), .ZN(new_n318));
  INV_X1    g0118(.A(G223), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n292), .B(new_n318), .C1(new_n319), .C2(new_n288), .ZN(new_n320));
  INV_X1    g0120(.A(new_n278), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G77), .C2(new_n292), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(new_n285), .C1(new_n214), .C2(new_n310), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n303), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n234), .B2(G50), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n326), .B2(new_n260), .C1(new_n262), .C2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n257), .B1(new_n213), .B2(new_n270), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n213), .B2(new_n267), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT68), .B(G179), .Z(new_n331));
  OAI211_X1 g0131(.A(new_n324), .B(new_n330), .C1(new_n323), .C2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n323), .A2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT9), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n334), .B1(new_n335), .B2(new_n323), .C1(new_n330), .C2(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n330), .A2(new_n336), .ZN(new_n338));
  OR3_X1    g0138(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT10), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n301), .A2(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n274), .C1(new_n335), .C2(new_n301), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G238), .A2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n292), .B(new_n344), .C1(new_n219), .C2(G1698), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G107), .B2(new_n292), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n321), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n284), .B1(new_n281), .B2(G244), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G200), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(G190), .A3(new_n350), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n267), .A2(new_n215), .ZN(new_n354));
  INV_X1    g0154(.A(new_n270), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G77), .ZN(new_n356));
  INV_X1    g0156(.A(new_n327), .ZN(new_n357));
  INV_X1    g0157(.A(new_n260), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n358), .B1(G20), .B2(G77), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT15), .B(G87), .Z(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n262), .B2(new_n361), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n354), .B(new_n356), .C1(new_n362), .C2(new_n257), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n352), .A2(new_n353), .A3(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n317), .A2(new_n341), .A3(new_n343), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n288), .A2(G226), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G33), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n367), .B(new_n368), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G87), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n259), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT73), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n373), .A2(new_n375), .ZN(new_n380));
  INV_X1    g0180(.A(new_n367), .ZN(new_n381));
  INV_X1    g0181(.A(new_n368), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  INV_X1    g0184(.A(new_n378), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n321), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n284), .B1(new_n281), .B2(G232), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(G190), .A3(new_n388), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n373), .A2(new_n258), .A3(new_n375), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n373), .A2(new_n394), .A3(new_n258), .A4(new_n375), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(G68), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n258), .B1(new_n234), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G159), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n260), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT72), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n397), .ZN(new_n402));
  OAI21_X1  g0202(.A(G20), .B1(new_n402), .B2(new_n233), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT72), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n399), .C2(new_n260), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  AND2_X1   g0208(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n409));
  NOR2_X1   g0209(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n259), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT3), .A2(G33), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(KEYINPUT7), .A3(new_n258), .A4(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n394), .B1(new_n292), .B2(G20), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n208), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n403), .B1(new_n399), .B2(new_n260), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n407), .A2(new_n257), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n267), .A2(new_n357), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n270), .B2(new_n357), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n390), .A2(new_n391), .A3(new_n418), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n366), .B1(new_n421), .B2(KEYINPUT74), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n391), .A2(new_n418), .A3(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT17), .A4(new_n390), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n363), .B1(new_n351), .B2(new_n303), .ZN(new_n427));
  INV_X1    g0227(.A(new_n331), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n349), .A2(new_n428), .A3(new_n350), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n387), .A2(new_n428), .A3(new_n388), .ZN(new_n431));
  AOI21_X1  g0231(.A(G169), .B1(new_n387), .B2(new_n388), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n418), .A2(new_n420), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT18), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n389), .A2(new_n303), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n387), .A2(new_n428), .A3(new_n388), .ZN(new_n437));
  AND4_X1   g0237(.A1(KEYINPUT18), .A2(new_n436), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n426), .B(new_n430), .C1(new_n435), .C2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n365), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n355), .B(new_n266), .C1(G1), .C2(new_n259), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT25), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n355), .B2(G107), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n442), .A2(G107), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(new_n283), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n278), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G264), .ZN(new_n455));
  INV_X1    g0255(.A(G257), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n373), .A2(new_n375), .B1(new_n456), .B2(G1698), .ZN(new_n457));
  OR2_X1    g0257(.A1(G250), .A2(G1698), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n457), .A2(new_n458), .B1(G33), .B2(G294), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n452), .B(new_n455), .C1(new_n459), .C2(new_n278), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n460), .A2(new_n335), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n377), .A2(G20), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n409), .A2(new_n410), .A3(new_n259), .ZN(new_n464));
  OAI211_X1 g0264(.A(KEYINPUT22), .B(new_n463), .C1(new_n464), .C2(new_n374), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n258), .A2(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT23), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n258), .A2(G33), .A3(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n292), .A2(new_n463), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT22), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT24), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT22), .B1(new_n292), .B2(new_n463), .ZN(new_n474));
  INV_X1    g0274(.A(new_n463), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n373), .B2(new_n375), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n476), .B2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n467), .A4(new_n468), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n462), .B1(new_n480), .B2(new_n257), .ZN(new_n481));
  AOI211_X1 g0281(.A(KEYINPUT79), .B(new_n266), .C1(new_n473), .C2(new_n479), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n446), .B(new_n461), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n460), .A2(G200), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n446), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n460), .A2(new_n303), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(G179), .B2(new_n460), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n209), .A2(new_n288), .ZN(new_n491));
  OAI221_X1 g0291(.A(new_n491), .B1(G244), .B2(new_n288), .C1(new_n464), .C2(new_n374), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n278), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n278), .B1(G250), .B2(new_n448), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n447), .A2(G1), .A3(G274), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(G200), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n441), .A2(new_n377), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(G20), .B(new_n208), .C1(new_n373), .C2(new_n375), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT19), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(new_n258), .A3(G33), .A4(G97), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(new_n377), .B1(new_n286), .B2(new_n258), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(new_n502), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n257), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n355), .A2(new_n360), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT76), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n258), .B(G68), .C1(new_n464), .C2(new_n374), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n266), .B1(new_n512), .B2(new_n506), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT76), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n513), .A2(new_n514), .A3(new_n509), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n498), .B(new_n500), .C1(new_n511), .C2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT77), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n497), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n492), .A2(new_n493), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n278), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n335), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n508), .A2(KEYINPUT76), .A3(new_n510), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n514), .B1(new_n513), .B2(new_n509), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n499), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(KEYINPUT77), .A3(new_n498), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n511), .A2(new_n515), .B1(new_n361), .B2(new_n441), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n428), .B(new_n519), .C1(new_n520), .C2(new_n278), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n303), .B1(new_n494), .B2(new_n497), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n530), .A2(KEYINPUT75), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT75), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n355), .A2(G97), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n358), .A2(G77), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n202), .A2(new_n203), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n504), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G20), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n413), .A2(new_n414), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n537), .B(new_n542), .C1(new_n543), .C2(new_n203), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n536), .B1(new_n544), .B2(new_n257), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n442), .A2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n288), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n216), .B1(new_n373), .B2(new_n375), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(KEYINPUT4), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n292), .B2(G250), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n553), .B2(new_n288), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n321), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n454), .A2(G257), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(new_n428), .A3(new_n452), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n452), .A3(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n303), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n547), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n555), .A2(G190), .A3(new_n452), .A4(new_n556), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n545), .A3(new_n546), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n453), .A2(new_n244), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n373), .A2(new_n375), .B1(new_n210), .B2(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n456), .A2(new_n288), .ZN(new_n568));
  INV_X1    g0368(.A(new_n292), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n567), .A2(new_n568), .B1(G303), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n452), .B(new_n566), .C1(new_n570), .C2(new_n278), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n270), .A2(G116), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n441), .B2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n256), .A2(new_n229), .B1(G20), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT78), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n551), .B(new_n258), .C1(G33), .C2(new_n202), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n576), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n577), .A2(new_n578), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n572), .B(new_n586), .C1(new_n335), .C2(new_n571), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(G169), .A3(new_n571), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G179), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n571), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n585), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n585), .A2(new_n571), .A3(KEYINPUT21), .A4(G169), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n587), .A2(new_n590), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n564), .A2(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n440), .A2(new_n490), .A3(new_n535), .A4(new_n596), .ZN(G372));
  INV_X1    g0397(.A(new_n430), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n343), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n317), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n317), .A2(KEYINPUT82), .A3(new_n599), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n426), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n435), .B2(new_n438), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n436), .A2(new_n434), .A3(new_n437), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT18), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n436), .A2(new_n434), .A3(KEYINPUT18), .A4(new_n437), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n339), .A2(new_n340), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n333), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n547), .A2(new_n557), .A3(new_n559), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n528), .A2(new_n534), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n486), .A2(new_n489), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n485), .A2(new_n484), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n622), .B2(new_n563), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n500), .B1(new_n511), .B2(new_n515), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT80), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n526), .A2(KEYINPUT80), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n523), .B(new_n498), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n616), .B(new_n619), .C1(new_n623), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n440), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n615), .A2(new_n632), .ZN(G369));
  NAND3_X1  g0433(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n269), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n229), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g0438(.A(G213), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n636), .B2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n586), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n595), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT84), .Z(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n480), .A2(new_n257), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT79), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n480), .A2(new_n462), .A3(new_n257), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n488), .B1(new_n655), .B2(new_n446), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n655), .A2(new_n446), .A3(new_n485), .A4(new_n461), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n486), .A2(new_n644), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n656), .B2(new_n645), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n645), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n634), .A2(new_n645), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n490), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n224), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR4_X1   g0469(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G1), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n235), .B2(new_n669), .ZN(new_n672));
  XOR2_X1   g0472(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n673));
  XNOR2_X1  g0473(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n619), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n657), .B(new_n563), .C1(new_n656), .C2(new_n634), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n560), .ZN(new_n677));
  INV_X1    g0477(.A(new_n630), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI211_X1 g0479(.A(KEYINPUT29), .B(new_n644), .C1(new_n679), .C2(new_n616), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT29), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n528), .A2(new_n534), .A3(new_n629), .A4(new_n617), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n624), .A2(new_n625), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n526), .A2(KEYINPUT80), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n522), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n560), .B1(new_n685), .B2(new_n498), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n616), .B(new_n682), .C1(new_n686), .C2(new_n629), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n628), .A2(new_n617), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT87), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n616), .A4(new_n682), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n628), .A2(new_n616), .ZN(new_n693));
  INV_X1    g0493(.A(new_n564), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n622), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n688), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n681), .B1(new_n696), .B2(new_n645), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n680), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  INV_X1    g0500(.A(new_n459), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n701), .A2(new_n321), .B1(G264), .B2(new_n454), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n592), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n494), .A2(new_n497), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n452), .A3(new_n556), .A4(new_n555), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n558), .A2(new_n521), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n592), .A3(KEYINPUT30), .A4(new_n702), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n460), .A2(new_n428), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n521), .A3(new_n558), .A4(new_n571), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n711), .A2(KEYINPUT86), .A3(new_n644), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT86), .B1(new_n711), .B2(new_n644), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT31), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n644), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT86), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(KEYINPUT86), .A3(new_n644), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n490), .A2(new_n535), .A3(new_n596), .A4(new_n645), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n714), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n699), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n674), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR3_X1   g0526(.A1(new_n269), .A2(new_n447), .A3(G20), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT88), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT88), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(G1), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n668), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n650), .B(new_n732), .C1(G330), .C2(new_n648), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT89), .Z(new_n734));
  OAI21_X1  g0534(.A(new_n230), .B1(new_n258), .B2(G169), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT90), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n428), .A2(new_n258), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT93), .Z(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n335), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n591), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(G326), .B1(G294), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT94), .Z(new_n745));
  NOR2_X1   g0545(.A1(new_n258), .A2(G179), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G329), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n745), .A2(new_n569), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n737), .A2(new_n747), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n737), .A2(new_n741), .ZN(new_n755));
  INV_X1    g0555(.A(G322), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n746), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT92), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT92), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n763), .A2(G303), .B1(G283), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n737), .A2(new_n765), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n751), .A2(new_n754), .A3(new_n757), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n738), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G50), .B1(G107), .B2(new_n770), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n569), .B1(new_n759), .B2(G87), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n208), .C2(new_n772), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n749), .A2(G159), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT91), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT32), .Z(new_n782));
  INV_X1    g0582(.A(new_n743), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n202), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n218), .A2(new_n755), .B1(new_n752), .B2(new_n215), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n779), .A2(new_n782), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n736), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n648), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(G355), .A2(new_n292), .A3(new_n224), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n254), .A2(new_n447), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n380), .A2(new_n667), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G45), .B2(new_n235), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(G116), .B2(new_n224), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n736), .A2(new_n790), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n787), .A2(new_n792), .A3(new_n731), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n734), .A2(new_n800), .ZN(G396));
  AOI21_X1  g0601(.A(new_n644), .B1(new_n679), .B2(new_n616), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n645), .A2(new_n363), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n353), .A2(new_n363), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n764), .B1(new_n349), .B2(new_n350), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n430), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT98), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n427), .A2(new_n429), .A3(new_n645), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n631), .A2(new_n645), .A3(new_n812), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n813), .A2(new_n724), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n732), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT100), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n813), .A2(new_n814), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n724), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n772), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n776), .A2(G303), .B1(new_n820), .B2(G283), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n575), .B2(new_n752), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT96), .Z(new_n823));
  AOI211_X1 g0623(.A(new_n292), .B(new_n823), .C1(G107), .C2(new_n763), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n753), .B2(new_n748), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n769), .A2(new_n377), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n755), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n825), .A2(new_n784), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n380), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n763), .B2(G50), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n770), .A2(G68), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n748), .ZN(new_n834));
  INV_X1    g0634(.A(new_n755), .ZN(new_n835));
  XOR2_X1   g0635(.A(KEYINPUT97), .B(G143), .Z(new_n836));
  AOI22_X1  g0636(.A1(new_n776), .A2(G137), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n326), .B2(new_n772), .C1(new_n399), .C2(new_n752), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  AOI211_X1 g0639(.A(new_n834), .B(new_n839), .C1(G58), .C2(new_n743), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n736), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n736), .A2(new_n788), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n215), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n810), .A2(new_n811), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n788), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n731), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n819), .A2(new_n847), .ZN(G384));
  NAND2_X1  g0648(.A1(new_n718), .A2(KEYINPUT101), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n711), .A2(new_n644), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n715), .A2(KEYINPUT101), .A3(new_n718), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n721), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n275), .A2(new_n644), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n317), .A2(new_n343), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n275), .B(new_n644), .C1(new_n307), .C2(new_n316), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n852), .A2(new_n812), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT81), .B1(new_n609), .B2(new_n610), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n610), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n426), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n642), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n434), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n642), .B1(new_n431), .B2(new_n432), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n434), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n421), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n421), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n407), .A2(new_n257), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n396), .B2(new_n406), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n420), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n422), .A2(new_n425), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n435), .A2(new_n438), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n861), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n863), .A2(new_n874), .B1(new_n423), .B2(new_n390), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n869), .B1(new_n878), .B2(new_n868), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n857), .B(KEYINPUT40), .C1(new_n871), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n877), .B2(new_n879), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n852), .A2(new_n812), .A3(new_n856), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n440), .A2(new_n852), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT102), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G330), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT103), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n440), .B1(new_n680), .B2(new_n697), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n615), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n317), .A2(new_n644), .ZN(new_n896));
  INV_X1    g0696(.A(new_n883), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n862), .A2(new_n870), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n896), .B(new_n899), .C1(new_n902), .C2(KEYINPUT39), .ZN(new_n903));
  INV_X1    g0703(.A(new_n884), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n644), .B(new_n844), .C1(new_n679), .C2(new_n616), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n427), .A2(new_n429), .A3(new_n645), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n904), .B(new_n856), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n612), .A2(new_n861), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n895), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n279), .B2(new_n635), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n575), .B1(new_n541), .B2(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n232), .C1(KEYINPUT35), .C2(new_n541), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n397), .A2(G77), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n235), .A2(new_n916), .B1(G50), .B2(new_n208), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n269), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n915), .A3(new_n918), .ZN(G367));
  XNOR2_X1  g0719(.A(new_n668), .B(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n665), .A2(new_n662), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n547), .A2(new_n644), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n694), .A2(new_n922), .B1(new_n617), .B2(new_n644), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT44), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n921), .A2(new_n923), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(new_n661), .Z(new_n929));
  OAI21_X1  g0729(.A(new_n665), .B1(new_n660), .B2(new_n664), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n650), .B(new_n930), .Z(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n698), .A3(new_n723), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(KEYINPUT104), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(KEYINPUT104), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n725), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n920), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n730), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n694), .A2(new_n922), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n665), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n560), .B1(new_n940), .B2(new_n620), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n645), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n683), .A2(new_n684), .A3(new_n644), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n693), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n616), .B2(new_n945), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n942), .A2(new_n944), .B1(KEYINPUT43), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n661), .A2(new_n923), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n950), .B(new_n951), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n939), .A2(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n213), .A2(new_n752), .B1(new_n772), .B2(new_n399), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT107), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n740), .A2(new_n836), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n770), .A2(G77), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n955), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n783), .A2(new_n208), .B1(new_n758), .B2(new_n218), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n569), .B(new_n960), .C1(new_n835), .C2(G150), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n956), .B(new_n962), .C1(G137), .C2(new_n749), .ZN(new_n963));
  INV_X1    g0763(.A(G317), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n830), .B1(new_n964), .B2(new_n748), .C1(new_n769), .C2(new_n202), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT106), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n739), .A2(new_n753), .ZN(new_n967));
  INV_X1    g0767(.A(G303), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n755), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  NOR4_X1   g0770(.A1(new_n966), .A2(new_n967), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n972));
  NAND2_X1  g0772(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n758), .C2(new_n575), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(new_n974), .C1(new_n827), .C2(new_n772), .ZN(new_n975));
  INV_X1    g0775(.A(new_n752), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(G283), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n743), .A2(G107), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n963), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n736), .ZN(new_n982));
  INV_X1    g0782(.A(new_n795), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n798), .B1(new_n224), .B2(new_n361), .C1(new_n245), .C2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n731), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n947), .A2(new_n791), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n953), .A2(new_n988), .ZN(G387));
  NAND2_X1  g0789(.A1(new_n743), .A2(new_n360), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n755), .B2(new_n213), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT109), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n380), .B1(new_n215), .B2(new_n758), .C1(new_n326), .C2(new_n748), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n976), .B2(G68), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n776), .A2(G159), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n820), .A2(new_n357), .B1(new_n770), .B2(G97), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n835), .A2(G317), .B1(new_n820), .B2(G311), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n968), .B2(new_n752), .C1(new_n739), .C2(new_n756), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n783), .C1(new_n827), .C2(new_n758), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n770), .A2(G116), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n749), .A2(G326), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n830), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n997), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n795), .B1(new_n241), .B2(new_n447), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n670), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1011), .A2(new_n224), .A3(new_n292), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n327), .A2(G50), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n447), .C1(new_n208), .C2(new_n215), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(G107), .B2(new_n224), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1009), .A2(new_n736), .B1(new_n798), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1019), .B(new_n731), .C1(new_n660), .C2(new_n791), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n931), .A2(new_n730), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n725), .A2(new_n931), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n668), .A3(new_n932), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(G393));
  NAND2_X1  g0825(.A1(new_n929), .A2(new_n932), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n933), .A2(new_n934), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n668), .B(new_n1026), .C1(new_n1027), .C2(new_n929), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n738), .A2(new_n964), .B1(new_n755), .B2(new_n753), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT52), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n770), .A2(G107), .B1(G322), .B2(new_n749), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n569), .A3(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n976), .A2(G294), .B1(G116), .B2(new_n743), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n968), .B2(new_n772), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT110), .Z(new_n1035));
  AOI211_X1 g0835(.A(new_n1032), .B(new_n1035), .C1(G283), .C2(new_n759), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n738), .A2(new_n326), .B1(new_n755), .B2(new_n399), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT51), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n820), .A2(G50), .B1(G68), .B2(new_n759), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n749), .A2(new_n836), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n215), .C2(new_n783), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n380), .B1(new_n752), .B2(new_n327), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n826), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1036), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT111), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n736), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n732), .B1(new_n923), .B2(new_n790), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n798), .B1(new_n202), .B2(new_n224), .C1(new_n251), .C2(new_n983), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n929), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n730), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1028), .A2(new_n1053), .ZN(G390));
  INV_X1    g0854(.A(new_n856), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n814), .B2(new_n809), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n865), .B(new_n642), .C1(new_n612), .C2(new_n426), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n870), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n901), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT39), .B1(new_n1059), .B2(new_n898), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT39), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n880), .A2(new_n883), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1056), .A2(new_n896), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n696), .A2(new_n645), .A3(new_n812), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n809), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n856), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n902), .A2(new_n896), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n852), .A2(new_n812), .A3(G330), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n856), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n440), .A2(G330), .A3(new_n852), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n893), .A2(new_n615), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1065), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT112), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n722), .A2(G330), .A3(new_n812), .A4(new_n856), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1070), .A2(new_n1055), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1055), .B1(new_n723), .B2(new_n844), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1071), .A2(new_n856), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n906), .B1(new_n802), .B2(new_n812), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1079), .A2(new_n1064), .A3(new_n1078), .A4(new_n809), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT112), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1063), .A2(new_n1068), .A3(new_n1078), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1072), .A2(new_n1075), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n896), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1084), .B2(new_n1055), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n899), .B1(new_n902), .B2(KEYINPUT39), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1093), .A2(new_n1094), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1095), .B2(new_n1082), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1089), .A2(new_n1075), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1098), .A3(new_n668), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT113), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n569), .B1(new_n976), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n758), .A2(new_n326), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT53), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n776), .A2(G128), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G132), .B2(new_n835), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n749), .A2(G125), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n770), .A2(G50), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n820), .A2(G137), .B1(G159), .B2(new_n743), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n820), .A2(G107), .B1(G77), .B2(new_n743), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1113), .B1(new_n377), .B2(new_n762), .C1(new_n575), .C2(new_n755), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n752), .A2(new_n202), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n738), .A2(new_n1001), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n832), .B(new_n569), .C1(new_n827), .C2(new_n748), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n736), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n865), .B1(new_n612), .B2(new_n426), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1058), .B1(new_n1120), .B2(new_n861), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n898), .B1(new_n1121), .B2(KEYINPUT38), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1062), .B1(new_n1122), .B2(new_n1061), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n731), .B(new_n1119), .C1(new_n1123), .C2(new_n789), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n842), .A2(new_n327), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1100), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1119), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1094), .B2(new_n788), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1129), .A2(KEYINPUT113), .A3(new_n731), .A4(new_n1125), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT114), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1090), .B(new_n730), .C1(new_n1095), .C2(new_n1082), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1099), .B1(new_n1134), .B2(new_n1135), .ZN(G378));
  OAI21_X1  g0936(.A(new_n1075), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n881), .A2(G330), .A3(new_n886), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n341), .B(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n330), .A2(new_n861), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1138), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1145), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n881), .A3(G330), .A4(new_n886), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(new_n910), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1137), .A2(new_n1150), .A3(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1146), .A2(new_n910), .A3(KEYINPUT118), .A4(new_n1148), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1091), .B2(new_n1075), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1151), .B(new_n668), .C1(new_n1156), .C2(KEYINPUT57), .ZN(new_n1157));
  AND4_X1   g0957(.A1(KEYINPUT118), .A2(new_n1146), .A3(new_n910), .A4(new_n1148), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1148), .A2(new_n1146), .B1(new_n910), .B2(KEYINPUT118), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n730), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n743), .A2(G68), .B1(new_n749), .B2(G283), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n277), .C1(new_n215), .C2(new_n758), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n755), .A2(new_n203), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT115), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n820), .A2(G97), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n770), .A2(G58), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n380), .B1(new_n776), .B2(G116), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1163), .B(new_n1169), .C1(new_n360), .C2(new_n976), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n213), .B1(new_n464), .B2(G41), .ZN(new_n1173));
  INV_X1    g0973(.A(G124), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n259), .B1(new_n748), .B2(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n835), .A2(G128), .B1(new_n976), .B2(G137), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n759), .A2(new_n1101), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n776), .A2(G125), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n820), .A2(G132), .B1(G150), .B2(new_n743), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G41), .B(new_n1175), .C1(new_n1180), .C2(KEYINPUT59), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(KEYINPUT59), .B2(new_n1180), .C1(new_n399), .C2(new_n769), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1172), .A2(new_n1173), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT117), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n736), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n842), .A2(new_n213), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1145), .A2(new_n788), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n731), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1157), .A2(new_n1161), .A3(new_n1188), .ZN(G375));
  NAND4_X1  g0989(.A1(new_n1074), .A2(new_n1086), .A3(new_n1080), .A4(new_n1088), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1097), .A2(new_n920), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n292), .B1(new_n776), .B2(G294), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n958), .C1(new_n968), .C2(new_n748), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n203), .A2(new_n752), .B1(new_n772), .B2(new_n575), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT120), .Z(new_n1195));
  OAI211_X1 g0995(.A(new_n1195), .B(new_n990), .C1(new_n202), .C2(new_n762), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(G283), .C2(new_n835), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT121), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1167), .B1(new_n213), .B2(new_n783), .C1(new_n833), .C2(new_n738), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G137), .B2(new_n835), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n820), .A2(new_n1101), .B1(G128), .B2(new_n749), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1200), .A2(new_n380), .A3(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n326), .B2(new_n752), .C1(new_n399), .C2(new_n762), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n732), .B1(new_n1204), .B2(new_n736), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n789), .B2(new_n856), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n208), .B2(new_n842), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n730), .B(KEYINPUT119), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1089), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1191), .A2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G375), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT123), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1099), .A2(new_n1133), .A3(new_n1131), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(KEYINPUT123), .B2(new_n1211), .ZN(new_n1215));
  INV_X1    g1015(.A(G390), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n953), .A2(new_n1216), .A3(new_n988), .ZN(new_n1217));
  OR2_X1    g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1217), .A2(G384), .A3(G381), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT122), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(KEYINPUT122), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1221), .B2(new_n1222), .ZN(G407));
  AOI21_X1  g1023(.A(new_n639), .B1(new_n1215), .B2(new_n643), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(G407), .ZN(G409));
  NAND2_X1  g1025(.A1(new_n643), .A2(G213), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1137), .A2(new_n1160), .A3(new_n920), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1188), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1150), .B2(new_n1208), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1137), .A2(new_n1160), .A3(KEYINPUT124), .A4(new_n920), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1213), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1157), .A2(G378), .A3(new_n1161), .A4(new_n1188), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1233), .B2(new_n1213), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1226), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT126), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n669), .B1(new_n1190), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1097), .C1(new_n1241), .C2(new_n1190), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G384), .A2(new_n1209), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1243), .B2(new_n1209), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1209), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n847), .A3(new_n819), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(KEYINPUT126), .A3(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G2897), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1226), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1249), .A2(new_n1244), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(G213), .A3(new_n643), .A4(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1239), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1251), .B(new_n1226), .C1(new_n1237), .C2(new_n1238), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1233), .A2(new_n1213), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1251), .A4(new_n1226), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1256), .A2(new_n1258), .A3(new_n1259), .A4(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n952), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n937), .B2(new_n938), .ZN(new_n1267));
  OAI21_X1  g1067(.A(G390), .B1(new_n1267), .B2(new_n987), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1217), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1218), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1217), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT127), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1265), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1257), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1257), .A2(new_n1280), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1259), .A4(new_n1256), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1278), .A2(new_n1283), .ZN(G405));
  AND2_X1   g1084(.A1(G375), .A2(new_n1213), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1236), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1254), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1251), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1279), .ZN(G402));
endmodule


