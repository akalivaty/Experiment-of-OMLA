//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G221), .B1(new_n189), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G143), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n198), .B(new_n201), .C1(new_n203), .C2(new_n196), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT75), .B1(new_n207), .B2(G104), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n207), .A3(G104), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n209), .A3(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n212), .B1(new_n219), .B2(G101), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT10), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n202), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n224), .A2(new_n225), .B1(new_n203), .B2(new_n227), .ZN(new_n228));
  NOR4_X1   g042(.A1(new_n202), .A2(KEYINPUT64), .A3(new_n223), .A4(new_n226), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n214), .A2(new_n218), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(new_n206), .A3(new_n213), .A4(new_n216), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n219), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(G137), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n240), .A2(new_n242), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n244), .A3(new_n242), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n246), .A2(new_n247), .B1(G131), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n205), .B2(new_n220), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n222), .A2(new_n237), .A3(new_n249), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(G131), .ZN(new_n253));
  INV_X1    g067(.A(new_n247), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n204), .B1(new_n232), .B2(new_n212), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT76), .B(new_n256), .C1(new_n221), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT77), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n261), .B(new_n256), .C1(new_n221), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n258), .B2(KEYINPUT77), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n266), .B(new_n268), .Z(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n222), .A2(new_n237), .A3(new_n251), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT78), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n222), .A2(new_n237), .A3(new_n273), .A4(new_n251), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n256), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n252), .A2(new_n269), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n265), .A2(new_n270), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n194), .B1(new_n279), .B2(G469), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n249), .B1(new_n272), .B2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n252), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n270), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n252), .A2(KEYINPUT79), .A3(new_n269), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n285), .B(new_n286), .C1(new_n263), .C2(new_n264), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n192), .A3(new_n193), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n191), .B1(new_n280), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n291));
  AND2_X1   g105(.A1(KEYINPUT66), .A2(G119), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT66), .A2(G119), .ZN(new_n293));
  OAI21_X1  g107(.A(G116), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(G116), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT2), .B(G113), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n294), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n234), .A2(new_n302), .A3(new_n236), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT80), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n234), .A2(new_n302), .A3(new_n305), .A4(new_n236), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(KEYINPUT5), .A3(new_n296), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT66), .B(G119), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G116), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(G113), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(new_n301), .A3(new_n232), .A4(new_n212), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT81), .ZN(new_n314));
  INV_X1    g128(.A(new_n220), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n301), .A4(new_n312), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G122), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n307), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n301), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT83), .B1(new_n321), .B2(new_n220), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n313), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n319), .B(KEYINPUT8), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n315), .A2(KEYINPUT83), .A3(new_n301), .A4(new_n312), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n230), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT7), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n204), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n267), .A2(G224), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n327), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n327), .B2(new_n330), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n334), .A2(new_n335), .A3(new_n328), .ZN(new_n336));
  OR3_X1    g150(.A1(new_n320), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n307), .A2(new_n318), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n319), .B(KEYINPUT82), .Z(new_n339));
  AOI21_X1  g153(.A(KEYINPUT6), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n307), .A2(new_n318), .A3(new_n319), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n314), .A2(new_n317), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n306), .B2(new_n304), .ZN(new_n343));
  INV_X1    g157(.A(new_n339), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(new_n345), .B2(KEYINPUT6), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n334), .A2(new_n335), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n193), .B(new_n337), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G210), .B1(G237), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n344), .B1(new_n307), .B2(new_n318), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT6), .B1(new_n320), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n343), .B2(new_n344), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n347), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n358), .A2(new_n193), .A3(new_n350), .A4(new_n337), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n291), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n348), .B1(new_n354), .B2(new_n356), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n320), .A2(new_n332), .A3(new_n336), .ZN(new_n362));
  NOR4_X1   g176(.A1(new_n361), .A2(G902), .A3(new_n362), .A4(new_n351), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT84), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n187), .B(new_n290), .C1(new_n360), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n309), .A2(G128), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n367), .A2(KEYINPUT72), .B1(G119), .B2(new_n199), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(KEYINPUT72), .B2(new_n367), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT24), .B(G110), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(KEYINPUT16), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n200), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n309), .A2(KEYINPUT73), .A3(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT73), .B1(new_n309), .B2(G128), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G110), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n375), .A2(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n374), .A2(new_n200), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT74), .B(G110), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n369), .A2(new_n371), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT22), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(G137), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n387), .B2(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT25), .B1(new_n403), .B2(G902), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(G234), .B2(new_n193), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT25), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n402), .A3(new_n407), .A4(new_n193), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n406), .A2(G902), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n402), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT71), .ZN(new_n413));
  NAND2_X1  g227(.A1(G472), .A2(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n256), .A2(new_n230), .ZN(new_n415));
  INV_X1    g229(.A(new_n244), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n239), .A2(G137), .ZN(new_n417));
  OAI21_X1  g231(.A(G131), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n204), .B(new_n418), .C1(new_n254), .C2(new_n255), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT70), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n422));
  INV_X1    g236(.A(new_n302), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n424), .A3(new_n419), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n302), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n423), .A3(new_n419), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT28), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G237), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT67), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G237), .ZN(new_n434));
  AOI21_X1  g248(.A(G953), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G210), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT26), .B(G101), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n439), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT69), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(KEYINPUT69), .A3(new_n441), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n430), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G472), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n202), .A2(new_n223), .A3(new_n226), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n225), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT64), .B1(new_n202), .B2(new_n223), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n419), .B(new_n448), .C1(new_n249), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n448), .B1(new_n415), .B2(new_n419), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n302), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n428), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n440), .A2(new_n441), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n426), .B2(new_n429), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n413), .B(new_n414), .C1(new_n447), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G472), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n430), .B2(new_n445), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n466), .B(new_n459), .C1(new_n461), .C2(new_n460), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n413), .B1(new_n467), .B2(new_n414), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n458), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n456), .A2(new_n428), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT31), .ZN(new_n472));
  INV_X1    g286(.A(new_n444), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(new_n442), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n429), .A3(new_n426), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n456), .A2(new_n476), .A3(new_n428), .A4(new_n470), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n465), .A3(new_n193), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(new_n481), .A3(new_n465), .A4(new_n193), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n412), .B1(new_n469), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n267), .A2(G952), .ZN(new_n485));
  INV_X1    g299(.A(G234), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n431), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(G902), .B(G953), .C1(new_n486), .C2(new_n431), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT95), .Z(new_n490));
  XOR2_X1   g304(.A(KEYINPUT21), .B(G898), .Z(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n432), .A2(new_n434), .ZN(new_n495));
  AND2_X1   g309(.A1(KEYINPUT85), .A2(G143), .ZN(new_n496));
  NOR2_X1   g310(.A1(KEYINPUT85), .A2(G143), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n495), .A2(new_n498), .A3(G214), .A4(new_n267), .ZN(new_n499));
  INV_X1    g313(.A(G214), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n500), .B(G953), .C1(new_n432), .C2(new_n434), .ZN(new_n501));
  INV_X1    g315(.A(new_n496), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n499), .B(G131), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n435), .A2(G214), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n496), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(KEYINPUT88), .A3(G131), .A4(new_n499), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT17), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n243), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(new_n508), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n376), .A3(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(G125), .B(G140), .Z(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G146), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n390), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT87), .ZN(new_n519));
  AND2_X1   g333(.A1(KEYINPUT18), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n507), .A2(KEYINPUT86), .A3(new_n499), .A4(new_n520), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G113), .B(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(G104), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT90), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n515), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n505), .A2(new_n508), .A3(new_n512), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n516), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND2_X1  g348(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n374), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n200), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(new_n389), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n525), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n527), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n529), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n494), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  AOI211_X1 g360(.A(KEYINPUT20), .B(new_n546), .C1(new_n529), .C2(new_n542), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n515), .A2(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n549), .B2(new_n529), .ZN(new_n550));
  INV_X1    g364(.A(G475), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n545), .A2(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT91), .ZN(new_n553));
  INV_X1    g367(.A(new_n529), .ZN(new_n554));
  INV_X1    g368(.A(new_n527), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n515), .B2(new_n525), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n193), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n559), .C1(new_n545), .C2(new_n547), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n493), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n197), .A2(G128), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT92), .B1(new_n199), .B2(G143), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n197), .A3(G128), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(new_n239), .ZN(new_n567));
  XNOR2_X1  g381(.A(G116), .B(G122), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT14), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G122), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G116), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n207), .B1(new_n572), .B2(KEYINPUT14), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n570), .A2(new_n573), .B1(new_n207), .B2(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G134), .B1(new_n562), .B2(KEYINPUT13), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n566), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n568), .B(new_n207), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n566), .A2(new_n578), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n189), .A2(new_n405), .A3(G953), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n577), .B2(new_n582), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n193), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  INV_X1    g402(.A(G478), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n577), .A2(new_n582), .ZN(new_n592));
  INV_X1    g406(.A(new_n583), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n594), .B2(new_n584), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n595), .A2(KEYINPUT94), .B1(KEYINPUT15), .B2(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(KEYINPUT94), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n561), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n366), .A2(new_n484), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n478), .A2(new_n193), .ZN(new_n602));
  NAND2_X1  g416(.A1(KEYINPUT96), .A2(G472), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n412), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n290), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT97), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n594), .B2(new_n584), .ZN(new_n610));
  OAI211_X1 g424(.A(G478), .B(new_n193), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT98), .B(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n587), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n553), .A2(new_n560), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n493), .ZN(new_n617));
  INV_X1    g431(.A(new_n187), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n352), .B2(new_n359), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n607), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n552), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n595), .B(KEYINPUT94), .C1(KEYINPUT15), .C2(new_n589), .ZN(new_n626));
  INV_X1    g440(.A(new_n597), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n590), .B1(new_n587), .B2(new_n588), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n493), .B(KEYINPUT99), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n619), .A2(new_n625), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n607), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n634), .B(new_n636), .ZN(G9));
  NAND2_X1  g451(.A1(new_n388), .A2(new_n396), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n401), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n410), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n409), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n366), .A2(new_n599), .A3(new_n604), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT101), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  XNOR2_X1  g460(.A(KEYINPUT102), .B(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n490), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n487), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n558), .B(new_n649), .C1(new_n545), .C2(new_n547), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n598), .A2(new_n650), .A3(KEYINPUT103), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n652));
  INV_X1    g466(.A(new_n649), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n552), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n654), .B2(new_n629), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n619), .A2(new_n642), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n469), .A2(new_n483), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n290), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n359), .A2(new_n291), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n357), .B2(new_n347), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n350), .B1(new_n663), .B2(new_n337), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n363), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n661), .B(new_n662), .C1(new_n665), .C2(new_n291), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n360), .B2(new_n364), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(KEYINPUT38), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT38), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n553), .A2(new_n560), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n649), .B(KEYINPUT39), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n290), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n670), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n642), .A2(new_n598), .ZN(new_n677));
  INV_X1    g491(.A(new_n457), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n427), .A2(new_n428), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n678), .A2(new_n470), .B1(new_n679), .B2(new_n474), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n680), .B2(G902), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n483), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n187), .A3(new_n677), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND4_X1  g498(.A1(new_n553), .A2(new_n560), .A3(new_n614), .A4(new_n649), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n657), .A2(new_n658), .A3(new_n290), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  AOI21_X1  g502(.A(new_n192), .B1(new_n288), .B2(new_n193), .ZN(new_n689));
  AOI211_X1 g503(.A(G469), .B(G902), .C1(new_n283), .C2(new_n287), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n690), .A3(new_n191), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n480), .A2(new_n482), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n414), .B1(new_n447), .B2(new_n462), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT71), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n463), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n605), .B(new_n691), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n620), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT41), .B(G113), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n632), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT105), .B(G116), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  OAI211_X1 g516(.A(new_n561), .B(new_n598), .C1(new_n692), .C2(new_n695), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n619), .A2(new_n642), .A3(new_n691), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n295), .ZN(G21));
  NAND4_X1  g520(.A1(new_n672), .A2(new_n619), .A3(new_n629), .A4(new_n631), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n602), .B(new_n465), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n605), .A3(new_n691), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n571), .ZN(G24));
  AND3_X1   g525(.A1(new_n619), .A2(new_n642), .A3(new_n691), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n712), .B(new_n708), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  OAI211_X1 g530(.A(new_n187), .B(new_n662), .C1(new_n665), .C2(new_n291), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n605), .B1(new_n692), .B2(new_n695), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n685), .B(KEYINPUT106), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(KEYINPUT42), .A3(new_n290), .A4(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n360), .A2(new_n364), .A3(new_n618), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n484), .A2(new_n723), .A3(new_n290), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n713), .A2(new_n714), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n290), .A3(new_n656), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  OR2_X1    g544(.A1(new_n279), .A2(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n279), .A2(KEYINPUT45), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(G469), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n194), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n690), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n191), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n673), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT107), .ZN(new_n741));
  INV_X1    g555(.A(new_n614), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n672), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT43), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n671), .A2(KEYINPUT43), .A3(new_n614), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n744), .A2(KEYINPUT108), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT108), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  INV_X1    g561(.A(new_n604), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n642), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n741), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n751), .A2(new_n717), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n241), .ZN(G39));
  OR2_X1    g568(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n658), .A2(new_n605), .A3(new_n685), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n723), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT109), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  OAI21_X1  g575(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n658), .A2(new_n598), .A3(new_n654), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n290), .A3(new_n642), .A4(new_n723), .ZN(new_n765));
  OAI22_X1  g579(.A1(new_n696), .A2(new_n632), .B1(new_n707), .B2(new_n709), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n697), .A3(new_n705), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n727), .A2(new_n765), .A3(new_n729), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n615), .B(KEYINPUT111), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n187), .B(new_n631), .C1(new_n360), .C2(new_n364), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n771), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n615), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT112), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n607), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n671), .A2(new_n629), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT113), .Z(new_n779));
  NAND3_X1  g593(.A1(new_n607), .A2(new_n779), .A3(new_n773), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n780), .A3(new_n600), .A4(new_n643), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n629), .B(new_n187), .C1(new_n664), .C2(new_n363), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n671), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n642), .A2(new_n653), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n290), .A3(new_n682), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n715), .A2(new_n786), .A3(new_n659), .A4(new_n687), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n768), .A2(new_n782), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n727), .A2(new_n765), .A3(new_n729), .A4(new_n767), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n781), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n789), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n789), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n792), .B2(new_n796), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(KEYINPUT116), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n804), .ZN(new_n809));
  INV_X1    g623(.A(new_n670), .ZN(new_n810));
  INV_X1    g624(.A(new_n709), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n488), .B(new_n811), .C1(new_n744), .C2(new_n745), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n618), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n813), .A4(new_n618), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n723), .A2(new_n691), .ZN(new_n819));
  INV_X1    g633(.A(new_n682), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n412), .A2(new_n487), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n819), .A2(KEYINPUT119), .A3(new_n820), .A4(new_n821), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n671), .A3(new_n742), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n744), .A2(new_n745), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n487), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n642), .A3(new_n708), .A4(new_n819), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n708), .A2(new_n605), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n827), .A2(new_n487), .A3(new_n831), .A4(new_n717), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n689), .A2(new_n690), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n191), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT118), .Z(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n757), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n818), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n824), .A2(new_n616), .A3(new_n825), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n755), .A2(new_n756), .A3(new_n835), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n842), .B2(new_n832), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n818), .A2(new_n843), .A3(new_n830), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n485), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n813), .A2(new_n619), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT120), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n828), .A2(new_n484), .A3(new_n819), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT48), .Z(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n806), .A2(new_n809), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT121), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n806), .A2(new_n809), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT122), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n412), .A2(new_n618), .A3(new_n191), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n682), .B1(new_n858), .B2(KEYINPUT110), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(KEYINPUT110), .B2(new_n858), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n833), .B(KEYINPUT49), .Z(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n810), .A2(new_n743), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n857), .A2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n357), .A2(new_n347), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n361), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT124), .Z(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n797), .A2(G902), .A3(new_n798), .ZN(new_n870));
  INV_X1    g684(.A(G210), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n872), .A2(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n873), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n867), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n267), .A2(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(G51));
  NAND2_X1  g696(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n808), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n288), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n870), .A2(new_n733), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n880), .B1(new_n888), .B2(new_n889), .ZN(G54));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n870), .A2(new_n891), .A3(new_n551), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n543), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n880), .ZN(G60));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n885), .A2(new_n808), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n608), .A2(new_n610), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(new_n881), .C1(new_n896), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n802), .B2(new_n884), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT125), .B1(new_n902), .B2(new_n880), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n806), .A2(new_n809), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n897), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n403), .B1(new_n799), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n909), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n797), .A2(new_n640), .A3(new_n798), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n881), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT126), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n910), .A2(new_n915), .A3(new_n881), .A4(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n914), .A2(KEYINPUT61), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(G66));
  AOI21_X1  g735(.A(new_n267), .B1(new_n491), .B2(G224), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n782), .A2(new_n767), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT127), .Z(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n924), .B2(new_n267), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n346), .B1(G898), .B2(new_n267), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(G69));
  NOR2_X1   g741(.A1(new_n454), .A2(new_n455), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n537), .Z(new_n929));
  INV_X1    g743(.A(new_n759), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n753), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n729), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n741), .A2(new_n484), .A3(new_n784), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n715), .A2(new_n659), .A3(new_n687), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n727), .A3(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n932), .A2(new_n935), .A3(G953), .ZN(new_n936));
  NAND2_X1  g750(.A1(G900), .A2(G953), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(G227), .A2(G900), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G953), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n674), .B(new_n719), .C1(new_n779), .C2(new_n775), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT62), .B1(new_n683), .B2(new_n934), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n683), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n931), .B(new_n942), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n267), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n939), .B(new_n941), .C1(new_n929), .C2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n932), .A2(new_n935), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n937), .B1(new_n948), .B2(G953), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(G953), .A3(new_n940), .A4(new_n929), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n947), .A2(new_n950), .ZN(G72));
  XOR2_X1   g765(.A(new_n414), .B(KEYINPUT63), .Z(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n945), .B2(new_n924), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n678), .A2(new_n458), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n952), .ZN(new_n956));
  AOI211_X1 g770(.A(new_n956), .B(new_n954), .C1(new_n792), .C2(new_n796), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n470), .B2(new_n457), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n881), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n952), .B1(new_n948), .B2(new_n924), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n457), .A2(new_n470), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(G57));
endmodule


