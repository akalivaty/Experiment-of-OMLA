//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n189), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n192), .B1(new_n201), .B2(new_n187), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n207), .B(G146), .C1(new_n203), .C2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n205), .A3(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n210), .A4(new_n211), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n202), .A2(KEYINPUT67), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n196), .B2(new_n200), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n188), .A2(G134), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n189), .B2(new_n198), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n197), .A2(KEYINPUT11), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n193), .B1(new_n195), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(new_n187), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT0), .A4(G128), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT65), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G113), .ZN(new_n238));
  INV_X1    g052(.A(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT2), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n231), .B(new_n233), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n224), .A2(new_n229), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n192), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n213), .A2(new_n223), .A3(new_n246), .A4(new_n216), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n217), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n217), .A2(new_n245), .A3(new_n249), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n256), .A2(new_n257), .A3(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n255), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n224), .B2(new_n229), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n217), .A2(new_n249), .A3(new_n264), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n196), .A2(new_n200), .A3(G131), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n187), .B1(new_n220), .B2(new_n222), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n229), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n212), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n214), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n223), .A3(new_n246), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n263), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n244), .A2(new_n236), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n265), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n254), .A2(new_n262), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT31), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n261), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n274), .B1(new_n268), .B2(new_n271), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT72), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n254), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n247), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT73), .B1(new_n268), .B2(new_n247), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(new_n275), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT28), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n265), .A2(new_n273), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n293), .A2(new_n275), .B1(new_n251), .B2(new_n253), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT31), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n262), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n277), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n280), .A2(new_n292), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n301), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n294), .B2(new_n262), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n282), .B1(new_n290), .B2(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n254), .A2(new_n286), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(KEYINPUT28), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n254), .A2(new_n276), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT29), .B1(new_n314), .B2(new_n261), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n316), .C1(new_n287), .C2(new_n310), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n217), .A2(new_n249), .A3(new_n268), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n275), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n254), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n291), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n261), .A2(new_n308), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n313), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n302), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n305), .A2(new_n307), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G478), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(KEYINPUT15), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(KEYINPUT15), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G902), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n232), .A2(KEYINPUT14), .A3(G122), .ZN(new_n335));
  XOR2_X1   g149(.A(G116), .B(G122), .Z(new_n336));
  OAI211_X1 g150(.A(G107), .B(new_n335), .C1(new_n336), .C2(KEYINPUT14), .ZN(new_n337));
  OR2_X1    g151(.A1(KEYINPUT82), .A2(G107), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT82), .A2(G107), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n207), .A2(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n203), .A2(G143), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(new_n190), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n190), .ZN(new_n345));
  OAI221_X1 g159(.A(new_n337), .B1(new_n336), .B2(new_n340), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n336), .B(new_n340), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT13), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n342), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n341), .A2(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(G134), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  INV_X1    g169(.A(G217), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n356), .A3(G953), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n346), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n346), .B2(new_n354), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n334), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT92), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n333), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n354), .ZN(new_n363));
  INV_X1    g177(.A(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n346), .A2(new_n354), .A3(new_n357), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n333), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT92), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n369), .A3(KEYINPUT93), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G475), .A2(G902), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT90), .Z(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT20), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n207), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G131), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n379), .B(G143), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n187), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT16), .ZN(new_n387));
  XNOR2_X1  g201(.A(G125), .B(G140), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n388), .A2(KEYINPUT19), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n388), .A2(KEYINPUT19), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n205), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT18), .A2(G131), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n388), .A2(new_n205), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n382), .A2(new_n395), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n382), .B2(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(G104), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n381), .A2(new_n383), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(KEYINPUT16), .B2(new_n386), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n205), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n380), .A2(KEYINPUT17), .A3(G131), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n390), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n406), .B(new_n402), .C1(new_n410), .C2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n378), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n406), .B1(new_n394), .B2(new_n402), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT89), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n376), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n408), .A2(new_n422), .A3(new_n416), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n417), .B1(new_n424), .B2(KEYINPUT20), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n402), .B1(new_n410), .B2(new_n415), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n426), .A2(new_n407), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n334), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G475), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G952), .ZN(new_n431));
  AOI211_X1 g245(.A(G953), .B(new_n431), .C1(G234), .C2(G237), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n334), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR4_X1   g249(.A1(new_n374), .A2(new_n425), .A3(new_n430), .A4(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n334), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n257), .A2(G227), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n338), .A3(new_n339), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT3), .B1(new_n405), .B2(G107), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n405), .C2(G107), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n444), .A2(new_n338), .A3(new_n452), .A4(new_n339), .ZN(new_n453));
  AOI21_X1  g267(.A(G101), .B1(new_n405), .B2(G107), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n446), .A2(new_n451), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(G104), .B1(new_n338), .B2(new_n339), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n405), .A2(G107), .ZN(new_n457));
  OAI21_X1  g271(.A(G101), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n214), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n204), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n269), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n270), .B1(new_n455), .B2(new_n458), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n224), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT12), .B(new_n224), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n455), .A2(new_n458), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n216), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT10), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n471), .A2(new_n472), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n224), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n405), .A2(G107), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n446), .A2(new_n451), .A3(new_n476), .A4(new_n453), .ZN(new_n477));
  INV_X1    g291(.A(G101), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n228), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n477), .A2(G101), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n470), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n443), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n475), .B1(new_n474), .B2(new_n483), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n443), .A2(new_n485), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n440), .B1(new_n491), .B2(G469), .ZN(new_n492));
  INV_X1    g306(.A(new_n484), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n443), .B1(new_n493), .B2(new_n489), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n484), .A2(KEYINPUT85), .A3(new_n486), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n470), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT85), .B1(new_n484), .B2(new_n486), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n439), .A3(new_n334), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n438), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n477), .A2(G101), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n455), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n274), .B1(new_n477), .B2(new_n479), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n455), .A2(new_n458), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT5), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(G113), .C1(KEYINPUT5), .C2(new_n231), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n241), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT86), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n510), .B1(new_n504), .B2(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n514), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n228), .A2(G125), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(G125), .B2(new_n270), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n257), .A2(G224), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT87), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n521), .B(new_n523), .Z(new_n524));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n512), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n514), .B(KEYINPUT8), .Z(new_n528));
  NAND2_X1  g342(.A1(new_n506), .A2(new_n509), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n511), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n520), .A2(KEYINPUT88), .B1(KEYINPUT7), .B2(new_n523), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(new_n521), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(G902), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G210), .B1(G237), .B2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n534), .A3(new_n536), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n436), .A2(new_n500), .A3(new_n501), .A4(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n230), .B2(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n230), .A2(G128), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  XNOR2_X1  g361(.A(G119), .B(G128), .ZN(new_n548));
  AOI22_X1  g362(.A1(G110), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n390), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n389), .A2(G146), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G110), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n543), .A2(new_n545), .A3(new_n553), .A4(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n554), .A2(new_n555), .B1(new_n547), .B2(new_n548), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n390), .B(new_n396), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(KEYINPUT77), .A3(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT22), .B(G137), .Z(new_n560));
  AND3_X1   g374(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT77), .B1(new_n552), .B2(new_n558), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(KEYINPUT77), .B(new_n563), .C1(new_n552), .C2(new_n558), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n334), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT25), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n565), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n559), .A3(new_n563), .ZN(new_n572));
  INV_X1    g386(.A(new_n567), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(KEYINPUT25), .A3(new_n334), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n356), .B1(G234), .B2(new_n334), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT80), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT79), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(G902), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT78), .Z(new_n582));
  AOI21_X1  g396(.A(new_n580), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n580), .A3(new_n582), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n578), .A2(new_n579), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  INV_X1    g401(.A(new_n577), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n570), .B2(new_n575), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT80), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n327), .A2(new_n541), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  NAND2_X1  g408(.A1(new_n298), .A2(new_n334), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n306), .ZN(new_n597));
  INV_X1    g411(.A(new_n500), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n597), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT94), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT95), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n538), .A2(new_n601), .A3(new_n539), .ZN(new_n602));
  INV_X1    g416(.A(new_n501), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n536), .B1(new_n527), .B2(new_n534), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n424), .A2(KEYINPUT20), .ZN(new_n607));
  INV_X1    g421(.A(new_n417), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n360), .A2(new_n328), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n365), .A2(new_n366), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT33), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(G478), .A3(new_n334), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n609), .A2(new_n429), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n606), .A2(new_n435), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND2_X1  g435(.A1(new_n420), .A2(new_n423), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n607), .B1(new_n622), .B2(new_n378), .ZN(new_n623));
  INV_X1    g437(.A(new_n435), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n374), .A3(new_n429), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n606), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n600), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n552), .A2(new_n558), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n582), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n578), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n634), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT97), .B1(new_n589), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n436), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n540), .A2(new_n501), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n598), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n298), .B2(new_n334), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n277), .A2(KEYINPUT31), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n311), .A2(KEYINPUT28), .ZN(new_n645));
  INV_X1    g459(.A(new_n291), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n647), .B2(new_n283), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n277), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT70), .B1(new_n277), .B2(KEYINPUT31), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n300), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n639), .A2(new_n641), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND3_X1  g470(.A1(new_n500), .A2(new_n635), .A3(new_n637), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT98), .B(G900), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n433), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n432), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n429), .A2(new_n623), .A3(new_n374), .A4(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n602), .A3(new_n605), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n327), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n302), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT75), .B1(new_n298), .B2(new_n302), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n301), .A2(new_n306), .B1(new_n324), .B2(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n657), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(KEYINPUT99), .A3(new_n664), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT100), .B(G128), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G30));
  INV_X1    g490(.A(new_n320), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n677), .A2(new_n678), .A3(new_n282), .ZN(new_n679));
  INV_X1    g493(.A(new_n277), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT101), .B1(new_n320), .B2(new_n283), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n682), .B2(G902), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n670), .A2(new_n307), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n578), .A2(new_n634), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n662), .B(KEYINPUT39), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n500), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n684), .B(new_n686), .C1(KEYINPUT40), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT38), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n540), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n538), .A2(KEYINPUT38), .A3(new_n539), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n425), .A2(new_n430), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n373), .B2(new_n372), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(new_n695), .A3(new_n501), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n207), .ZN(G45));
  INV_X1    g514(.A(new_n662), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n606), .A2(new_n617), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n672), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NAND2_X1  g518(.A1(new_n499), .A2(new_n437), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n498), .A2(new_n334), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(G469), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT102), .B(new_n439), .C1(new_n498), .C2(new_n334), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n705), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n327), .A2(new_n618), .A3(new_n592), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n327), .A2(new_n592), .A3(new_n626), .A4(new_n712), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT103), .B(G116), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G18));
  AND2_X1   g532(.A1(new_n499), .A2(new_n437), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n708), .B2(new_n710), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n606), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n327), .A2(new_n721), .A3(new_n639), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  OAI211_X1 g537(.A(new_n719), .B(new_n624), .C1(new_n708), .C2(new_n710), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n697), .A2(new_n602), .A3(new_n605), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n587), .A2(new_n589), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n321), .A2(new_n282), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n296), .A2(new_n278), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n299), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n643), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND3_X1  g548(.A1(new_n596), .A2(new_n685), .A3(new_n730), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n720), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n702), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  AOI21_X1  g552(.A(KEYINPUT32), .B1(new_n298), .B2(new_n299), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n303), .B1(new_n739), .B2(KEYINPUT104), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n741), .B(KEYINPUT32), .C1(new_n298), .C2(new_n299), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n652), .B2(KEYINPUT32), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(KEYINPUT104), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n303), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n325), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n616), .A2(new_n662), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n538), .A2(new_n501), .A3(new_n539), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n598), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(KEYINPUT42), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n748), .A2(new_n727), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n591), .B1(new_n670), .B2(new_n671), .ZN(new_n754));
  INV_X1    g568(.A(new_n749), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n598), .A2(new_n750), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND4_X1  g575(.A1(new_n327), .A2(new_n592), .A3(new_n663), .A4(new_n756), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  NAND2_X1  g577(.A1(new_n485), .A2(new_n443), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n489), .B2(new_n487), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n439), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n491), .A2(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n440), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n440), .B1(new_n767), .B2(new_n768), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n499), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n437), .A3(new_n687), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n696), .B2(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n612), .A2(new_n615), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n696), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n696), .B(new_n780), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n597), .A3(new_n685), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n597), .A3(KEYINPUT44), .A4(new_n685), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT107), .ZN(new_n789));
  INV_X1    g603(.A(new_n750), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n789), .B1(new_n788), .B2(new_n790), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n778), .B(new_n787), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  INV_X1    g610(.A(new_n775), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n499), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n796), .B1(new_n799), .B2(new_n438), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n437), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n591), .A2(new_n755), .A3(new_n790), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n327), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(new_n684), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n499), .B1(new_n708), .B2(new_n710), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n781), .A2(new_n603), .A3(new_n438), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n693), .A2(new_n727), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n713), .A2(new_n716), .A3(new_n722), .A4(new_n733), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n638), .B1(new_n670), .B2(new_n671), .ZN(new_n818));
  AOI21_X1  g632(.A(G902), .B1(new_n648), .B2(new_n651), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n727), .B(new_n730), .C1(new_n819), .C2(new_n642), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n697), .A2(new_n602), .A3(new_n605), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n818), .A2(new_n721), .B1(new_n822), .B2(new_n725), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n713), .A4(new_n716), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n751), .A2(new_n685), .A3(new_n732), .ZN(new_n826));
  INV_X1    g640(.A(new_n370), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n429), .A2(new_n623), .A3(new_n827), .A4(new_n662), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n637), .A3(new_n635), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n327), .A2(new_n756), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n762), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n425), .A2(new_n430), .A3(new_n827), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n624), .B1(new_n616), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n640), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n592), .A3(new_n500), .A4(new_n653), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n593), .A2(new_n835), .A3(new_n654), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n760), .A2(new_n817), .A3(new_n825), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n702), .B1(new_n672), .B2(new_n736), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n821), .A2(new_n598), .A3(new_n701), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n684), .A3(new_n686), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT99), .B1(new_n672), .B2(new_n664), .ZN(new_n842));
  AND4_X1   g656(.A1(KEYINPUT99), .A2(new_n327), .A3(new_n658), .A4(new_n664), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n839), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n674), .A2(KEYINPUT52), .A3(new_n839), .A4(new_n841), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT53), .B1(new_n838), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n816), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n760), .A3(new_n837), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n846), .B2(new_n847), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n849), .A2(new_n853), .A3(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n838), .A2(new_n848), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT110), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n857), .A3(new_n850), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n838), .B(new_n848), .C1(new_n856), .C2(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n854), .B1(new_n860), .B2(KEYINPUT54), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n750), .A2(new_n661), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n784), .A2(new_n712), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n727), .A3(new_n748), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n735), .B1(new_n864), .B2(new_n865), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n592), .A2(new_n809), .A3(new_n712), .A4(new_n862), .ZN(new_n870));
  INV_X1    g684(.A(new_n696), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n780), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT114), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n784), .A2(new_n732), .A3(new_n727), .A4(new_n432), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n694), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n712), .A2(KEYINPUT113), .A3(new_n603), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n720), .B2(new_n501), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n877), .A2(new_n875), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n876), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n810), .A2(new_n437), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n790), .B(new_n886), .C1(new_n802), .C2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n873), .A2(new_n885), .A3(KEYINPUT51), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n870), .A2(new_n616), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n431), .B(G953), .C1(new_n886), .C2(new_n721), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n868), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n894));
  INV_X1    g708(.A(new_n884), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n873), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n886), .A2(new_n790), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n887), .B1(new_n802), .B2(KEYINPUT112), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n893), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT117), .B(new_n893), .C1(new_n898), .C2(new_n902), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n892), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n861), .A2(new_n907), .A3(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n431), .A2(new_n257), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT118), .B1(new_n861), .B2(new_n907), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n815), .B1(new_n910), .B2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n257), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(G210), .B(G902), .C1(new_n849), .C2(new_n853), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n519), .A2(new_n526), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n524), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT120), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n920), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n917), .A2(KEYINPUT119), .A3(new_n920), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G51));
  NOR2_X1   g741(.A1(new_n849), .A2(new_n853), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT54), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n440), .B(KEYINPUT57), .Z(new_n930));
  OAI21_X1  g744(.A(new_n498), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n928), .A2(new_n334), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n768), .A3(new_n767), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n913), .B1(new_n931), .B2(new_n933), .ZN(G54));
  NAND3_X1  g748(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n622), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n622), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n913), .ZN(G60));
  XNOR2_X1  g752(.A(new_n614), .B(KEYINPUT121), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n914), .B1(new_n929), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(new_n854), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n939), .B2(new_n946), .ZN(G63));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT60), .Z(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n849), .B2(new_n853), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n952));
  INV_X1    g766(.A(new_n574), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n950), .C1(new_n849), .C2(new_n853), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n914), .ZN(new_n957));
  INV_X1    g771(.A(new_n633), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n952), .B2(new_n955), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n948), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n952), .A2(new_n955), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n633), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n914), .A4(new_n956), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(G66));
  INV_X1    g778(.A(new_n434), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n257), .B1(new_n965), .B2(G224), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n817), .A2(new_n825), .ZN(new_n967));
  INV_X1    g781(.A(new_n836), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(new_n257), .ZN(new_n971));
  INV_X1    g785(.A(G898), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n918), .B1(new_n972), .B2(G953), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n674), .A2(new_n839), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n674), .A2(KEYINPUT123), .A3(new_n839), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n760), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n778), .A2(new_n748), .A3(new_n727), .A4(new_n726), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n807), .A2(new_n794), .A3(new_n762), .A4(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT126), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n762), .A2(new_n807), .A3(new_n794), .A4(new_n982), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n980), .A3(new_n986), .A4(new_n760), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n987), .A3(new_n257), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n391), .A2(new_n392), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n293), .B(new_n989), .Z(new_n990));
  INV_X1    g804(.A(G900), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n257), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n975), .B1(new_n994), .B2(KEYINPUT125), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n616), .A2(new_n832), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n750), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n997), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(new_n688), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n754), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n807), .A2(new_n794), .A3(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n689), .A2(new_n698), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n980), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1004), .B2(KEYINPUT62), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n980), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n994), .B1(new_n1008), .B2(new_n990), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n995), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g824(.A(new_n994), .B1(KEYINPUT125), .B2(new_n975), .C1(new_n1008), .C2(new_n990), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1010), .A2(new_n1011), .ZN(G72));
  NAND3_X1  g826(.A1(new_n1005), .A2(new_n969), .A3(new_n1007), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n262), .A3(new_n314), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n294), .A2(new_n262), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n860), .B(new_n1015), .C1(new_n680), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n984), .A2(new_n987), .A3(new_n969), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1021), .A2(new_n1015), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n314), .A2(new_n262), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(KEYINPUT127), .B(new_n914), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n913), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n1025), .B2(new_n1028), .ZN(G57));
endmodule


