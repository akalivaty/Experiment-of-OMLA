//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT0), .A4(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n187), .A2(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT64), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n205), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT65), .B1(new_n207), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n197), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n222));
  OAI211_X1 g036(.A(G128), .B(new_n222), .C1(new_n192), .C2(new_n193), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(G134), .B2(new_n201), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n204), .A2(new_n229), .B1(new_n203), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n211), .A2(new_n221), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n207), .A2(new_n208), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n238), .A2(new_n196), .B1(new_n226), .B2(new_n231), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n220), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n211), .A2(KEYINPUT28), .A3(new_n221), .A4(new_n234), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G237), .A2(G953), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G210), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n211), .A2(KEYINPUT30), .A3(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n239), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n220), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT31), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n235), .A4(new_n247), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n235), .A3(new_n247), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n253), .A2(new_n259), .A3(new_n235), .A4(new_n247), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G472), .A2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(KEYINPUT32), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n253), .A2(new_n235), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n248), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n237), .A2(new_n247), .A3(new_n240), .A4(new_n241), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n274), .A3(new_n248), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n270), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n207), .A2(new_n208), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n208), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n196), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n233), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT66), .B1(new_n223), .B2(new_n225), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n284), .A3(new_n231), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n282), .A2(new_n285), .A3(new_n220), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n221), .B1(new_n211), .B2(new_n234), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n277), .B(KEYINPUT28), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n237), .A2(KEYINPUT69), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n220), .B1(new_n282), .B2(new_n285), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n236), .B1(new_n290), .B2(new_n235), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n248), .A2(new_n272), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n276), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT70), .B1(new_n295), .B2(G472), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  INV_X1    g111(.A(G472), .ZN(new_n298));
  AOI211_X1 g112(.A(new_n297), .B(new_n298), .C1(new_n276), .C2(new_n294), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n266), .B(new_n267), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT16), .ZN(new_n302));
  AND2_X1   g116(.A1(KEYINPUT71), .A2(G125), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT71), .A2(G125), .ZN(new_n304));
  OAI21_X1  g118(.A(G140), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OR2_X1    g119(.A1(G125), .A2(G140), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT71), .A2(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT71), .A2(G125), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT16), .B(G140), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n187), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n309), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n302), .A3(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G125), .A2(G140), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n312), .B2(G140), .ZN(new_n316));
  OAI211_X1 g130(.A(G146), .B(new_n314), .C1(new_n316), .C2(new_n302), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n212), .A2(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n224), .A2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT24), .B(G110), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n212), .B2(G128), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n319), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n323), .B1(G110), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g143(.A1(G125), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n331), .B2(new_n315), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n306), .A2(KEYINPUT72), .A3(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(G110), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n325), .A2(new_n326), .A3(new_n336), .A4(new_n319), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n334), .A2(new_n187), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n317), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n318), .A2(new_n328), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n317), .A2(new_n338), .A3(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G953), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT74), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G137), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n305), .A2(new_n306), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT16), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n352), .B2(new_n314), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n307), .A2(new_n310), .A3(new_n187), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n328), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n331), .A2(new_n315), .A3(new_n329), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT72), .B1(new_n306), .B2(new_n330), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n187), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n335), .A2(new_n337), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n340), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n355), .A2(new_n361), .A3(new_n342), .A4(new_n348), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n301), .B(new_n350), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n341), .A2(new_n368), .A3(new_n342), .A4(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n366), .A2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n343), .B2(new_n349), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n301), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT77), .B1(new_n379), .B2(new_n381), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n371), .A2(new_n350), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n381), .A2(G902), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT78), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n382), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  OAI21_X1  g203(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT79), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n394), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n228), .A2(new_n233), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT10), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n226), .A2(new_n405), .A3(KEYINPUT10), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT80), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n395), .A2(new_n398), .A3(new_n415), .A4(new_n400), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n413), .A2(new_n414), .A3(G101), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n399), .B1(new_n412), .B2(KEYINPUT80), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n420), .A2(KEYINPUT81), .A3(new_n414), .A4(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n420), .B2(new_n416), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n196), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n209), .A2(new_n210), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n411), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n411), .B2(new_n426), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n344), .A2(G227), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n226), .B(new_n405), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n278), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT12), .B1(new_n280), .B2(new_n281), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n437), .A2(KEYINPUT12), .B1(new_n438), .B2(new_n436), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n428), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT82), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n439), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n433), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n411), .A2(new_n426), .ZN(new_n444));
  INV_X1    g258(.A(new_n427), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n428), .A3(new_n435), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n393), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n435), .B1(new_n446), .B2(new_n428), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n428), .A2(new_n435), .A3(new_n439), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n393), .B(new_n301), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n393), .A2(new_n301), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n392), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G475), .ZN(new_n459));
  INV_X1    g273(.A(new_n318), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n461));
  INV_X1    g275(.A(G237), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n344), .A3(G214), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n189), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n243), .A2(G143), .A3(G214), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n466), .B2(G131), .ZN(new_n467));
  AOI211_X1 g281(.A(KEYINPUT89), .B(new_n229), .C1(new_n464), .C2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT17), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n465), .ZN(new_n470));
  AOI21_X1  g284(.A(G143), .B1(new_n243), .B2(G214), .ZN(new_n471));
  OAI21_X1  g285(.A(G131), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT89), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n229), .A3(new_n465), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n466), .A2(new_n461), .A3(G131), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n464), .A2(KEYINPUT88), .A3(new_n229), .A4(new_n465), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n473), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n460), .B(new_n469), .C1(KEYINPUT17), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(G146), .B1(new_n332), .B2(new_n333), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(G146), .B2(new_n316), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n466), .A2(KEYINPUT18), .A3(G131), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT18), .A2(G131), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n464), .A2(new_n465), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT87), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n358), .B1(new_n351), .B2(new_n187), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n485), .A4(new_n483), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G113), .B(G122), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n394), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n480), .A2(new_n494), .A3(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n459), .B1(new_n498), .B2(new_n301), .ZN(new_n499));
  INV_X1    g313(.A(new_n497), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n479), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n476), .A2(new_n478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n467), .A2(new_n468), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT90), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n316), .A2(KEYINPUT19), .ZN(new_n506));
  INV_X1    g320(.A(new_n334), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n187), .C1(new_n507), .C2(KEYINPUT19), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(new_n505), .A3(new_n317), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n494), .B1(new_n509), .B2(new_n491), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT20), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n317), .B(new_n508), .C1(new_n479), .C2(new_n501), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT90), .B1(new_n503), .B2(new_n504), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n491), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n495), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n497), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n512), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n499), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT95), .ZN(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(G952), .A3(new_n344), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT94), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n533));
  INV_X1    g347(.A(G122), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G116), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n214), .A2(G122), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n397), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n536), .A3(new_n397), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT91), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n541));
  INV_X1    g355(.A(new_n539), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n224), .A2(G143), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n199), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G128), .B(G143), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n214), .A2(KEYINPUT14), .A3(G122), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n535), .A2(new_n536), .ZN(new_n554));
  OAI211_X1 g368(.A(G107), .B(new_n553), .C1(new_n554), .C2(KEYINPUT14), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n548), .A2(G134), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n548), .A2(G134), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n539), .A4(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n389), .A2(new_n380), .A3(G953), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n540), .A2(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n562));
  INV_X1    g376(.A(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n533), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(KEYINPUT92), .B(G902), .C1(new_n560), .C2(new_n564), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n532), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n564), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n301), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT92), .B1(new_n571), .B2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g386(.A(new_n532), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n522), .A2(new_n530), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n458), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G210), .B1(G237), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n196), .A2(new_n312), .ZN(new_n581));
  INV_X1    g395(.A(new_n226), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n312), .ZN(new_n583));
  INV_X1    g397(.A(G224), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G953), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n583), .B(new_n585), .Z(new_n586));
  NOR2_X1   g400(.A1(new_n424), .A2(new_n221), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n422), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n212), .A3(G116), .ZN(new_n590));
  OAI211_X1 g404(.A(G113), .B(new_n590), .C1(new_n216), .C2(new_n589), .ZN(new_n591));
  AND4_X1   g405(.A1(new_n218), .A2(new_n591), .A3(new_n401), .A4(new_n404), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G122), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n588), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT84), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n588), .A2(new_n593), .ZN(new_n599));
  INV_X1    g413(.A(new_n594), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n592), .B1(new_n422), .B2(new_n587), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n597), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n586), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n594), .B(KEYINPUT8), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n218), .A2(new_n591), .B1(new_n401), .B2(new_n404), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n607), .B1(new_n592), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(KEYINPUT85), .B(new_n607), .C1(new_n592), .C2(new_n608), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT7), .B1(new_n584), .B2(G953), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n583), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT7), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n583), .B1(new_n615), .B2(new_n585), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(new_n612), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n592), .B(new_n600), .C1(new_n422), .C2(new_n587), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n301), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n580), .B1(new_n606), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n586), .ZN(new_n621));
  INV_X1    g435(.A(new_n597), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n603), .B2(new_n594), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n604), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n603), .A2(new_n594), .A3(new_n622), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n619), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n579), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n606), .A2(new_n619), .A3(new_n580), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT86), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(G214), .B1(G237), .B2(G902), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT83), .Z(new_n634));
  AND3_X1   g448(.A1(new_n629), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n300), .A2(new_n388), .A3(new_n578), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  INV_X1    g451(.A(new_n388), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n256), .B2(new_n261), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n298), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n262), .B2(new_n263), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n579), .B1(new_n626), .B2(new_n627), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n633), .B1(new_n630), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n458), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n494), .B1(new_n480), .B2(new_n491), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n301), .B1(new_n500), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(G475), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n520), .B1(new_n519), .B2(new_n512), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT20), .B(new_n513), .C1(new_n518), .C2(new_n497), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n564), .B2(KEYINPUT96), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n570), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n531), .A2(G902), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT97), .B(G478), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n571), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n529), .B2(new_n527), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n643), .A2(new_n646), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT98), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT34), .B(G104), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  OAI211_X1 g480(.A(new_n575), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n530), .B(KEYINPUT99), .Z(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n643), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NAND2_X1  g487(.A1(new_n379), .A2(new_n381), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT77), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n379), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n343), .B1(KEYINPUT36), .B2(new_n349), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n362), .A2(KEYINPUT36), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n386), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n676), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n578), .A2(new_n641), .A3(new_n682), .A4(new_n635), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n526), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n529), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n667), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n300), .A2(new_n646), .A3(new_n682), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  AND3_X1   g505(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n448), .B1(new_n443), .B2(new_n447), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n695), .B2(new_n452), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n455), .B1(new_n696), .B2(new_n393), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n391), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n688), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  INV_X1    g515(.A(new_n633), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n652), .A2(new_n575), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n682), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n258), .A2(new_n260), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n247), .B1(new_n290), .B2(new_n235), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n301), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G472), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n266), .A2(new_n267), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT100), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n629), .A2(new_n632), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT38), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT38), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n706), .A2(new_n712), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n189), .ZN(G45));
  INV_X1    g532(.A(new_n688), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n652), .A2(new_n660), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n300), .A2(new_n646), .A3(new_n682), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  OAI21_X1  g537(.A(new_n301), .B1(new_n451), .B2(new_n453), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n392), .A3(new_n454), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n645), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n300), .A2(new_n388), .A3(new_n662), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND4_X1  g544(.A1(new_n300), .A2(new_n388), .A3(new_n670), .A4(new_n727), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  INV_X1    g546(.A(new_n577), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n300), .A2(new_n733), .A3(new_n682), .A4(new_n727), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  OAI211_X1 g549(.A(new_n288), .B(new_n248), .C1(new_n289), .C2(new_n291), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n261), .A2(new_n255), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT101), .A3(new_n263), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT101), .B1(new_n737), .B2(new_n263), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n640), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n645), .A2(new_n703), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n726), .A2(new_n669), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n388), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT102), .B(G122), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G24));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n682), .A3(new_n721), .A4(new_n727), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT103), .B(G125), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G27));
  OAI21_X1  g563(.A(KEYINPUT104), .B1(new_n434), .B2(new_n440), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n447), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(G469), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n391), .B1(new_n697), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n713), .A2(new_n633), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n300), .A3(new_n388), .A4(new_n721), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n295), .A2(G472), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n297), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n295), .A2(KEYINPUT70), .A3(G472), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n267), .A2(KEYINPUT105), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n267), .A2(KEYINPUT105), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n266), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n702), .B1(new_n629), .B2(new_n632), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n721), .A3(new_n754), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n767), .A3(KEYINPUT42), .A4(new_n388), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND4_X1  g584(.A1(new_n755), .A2(new_n300), .A3(new_n388), .A4(new_n689), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  INV_X1    g586(.A(new_n660), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n652), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT43), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n642), .A4(new_n682), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n766), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT107), .B1(new_n776), .B2(new_n766), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n522), .A2(new_n660), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n681), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n382), .A2(new_n383), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n641), .A3(new_n784), .ZN(new_n785));
  OAI22_X1  g599(.A1(new_n777), .A2(new_n778), .B1(KEYINPUT44), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n750), .A2(KEYINPUT45), .A3(new_n752), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n441), .A2(new_n788), .A3(new_n449), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n789), .A3(G469), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(new_n787), .A3(KEYINPUT106), .A4(G469), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n455), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(KEYINPUT46), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n454), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n392), .B(new_n699), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n786), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n201), .ZN(G39));
  INV_X1    g613(.A(new_n300), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n638), .A3(new_n721), .A4(new_n766), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n392), .B1(new_n795), .B2(new_n796), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT47), .B(new_n392), .C1(new_n795), .C2(new_n796), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n313), .ZN(G42));
  NAND3_X1  g621(.A1(new_n774), .A2(new_n634), .A3(new_n392), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n725), .A2(new_n454), .ZN(new_n809));
  AOI211_X1 g623(.A(new_n808), .B(new_n638), .C1(KEYINPUT49), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT108), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n712), .A3(new_n716), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n529), .ZN(new_n814));
  INV_X1    g628(.A(new_n726), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n766), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n782), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n765), .A2(new_n388), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT48), .Z(new_n820));
  NOR2_X1   g634(.A1(new_n782), .A2(new_n529), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n741), .A2(new_n388), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n645), .A3(new_n726), .ZN(new_n824));
  INV_X1    g638(.A(G952), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n824), .A2(new_n825), .A3(G953), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n638), .A2(new_n816), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n712), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n820), .B(new_n826), .C1(new_n661), .C2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n809), .A2(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n809), .A2(KEYINPUT111), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n391), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n804), .A2(new_n805), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n822), .A3(new_n766), .A4(new_n821), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n633), .B1(KEYINPUT112), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n716), .A2(new_n815), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n822), .A3(new_n821), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n716), .A2(new_n815), .A3(new_n836), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n823), .A2(new_n840), .B1(KEYINPUT112), .B2(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n741), .A2(new_n682), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n817), .A2(KEYINPUT113), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT113), .B1(new_n817), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n827), .A2(new_n712), .A3(new_n522), .A4(new_n773), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n834), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n834), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n829), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n391), .B(new_n688), .C1(new_n697), .C2(new_n753), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n784), .A2(new_n742), .A3(new_n711), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n690), .A2(new_n722), .A3(new_n747), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n702), .B1(new_n620), .B2(new_n628), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n698), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n266), .A2(new_n267), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n762), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n682), .A2(new_n689), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n382), .A2(new_n383), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n720), .B1(new_n863), .B2(new_n681), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n747), .A4(new_n855), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n857), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n636), .A2(new_n728), .A3(new_n731), .A4(new_n683), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n667), .B1(new_n522), .B2(new_n773), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(new_n698), .A3(new_n668), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n388), .A3(new_n635), .A4(new_n641), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n873), .A2(new_n734), .A3(new_n744), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n755), .A2(new_n682), .A3(new_n721), .A4(new_n741), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n522), .A2(new_n576), .A3(new_n719), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n458), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n300), .A2(new_n878), .A3(new_n682), .A4(new_n766), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n771), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n758), .B2(new_n768), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n868), .A2(new_n869), .A3(new_n875), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n771), .A2(new_n876), .A3(new_n879), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n769), .A2(new_n883), .A3(new_n870), .A4(new_n874), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n857), .A2(new_n867), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT53), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n869), .A2(KEYINPUT109), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n882), .A2(new_n886), .B1(new_n868), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n868), .A2(new_n884), .A3(KEYINPUT109), .A4(new_n869), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n882), .B2(new_n886), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n853), .A2(new_n891), .A3(KEYINPUT114), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n825), .A2(new_n344), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n890), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n894), .B1(new_n900), .B2(KEYINPUT54), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT114), .B1(new_n901), .B2(new_n853), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n813), .B1(new_n898), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n344), .A2(G952), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n882), .A2(new_n886), .A3(G902), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n882), .A2(new_n886), .A3(new_n907), .A4(G902), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n580), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n625), .B1(new_n601), .B2(new_n598), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n586), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n626), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n882), .A2(new_n886), .A3(G210), .A4(G902), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(KEYINPUT115), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n916), .B2(KEYINPUT115), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n915), .A2(KEYINPUT117), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G51));
  XNOR2_X1  g739(.A(new_n455), .B(KEYINPUT57), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n882), .A2(new_n886), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n892), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n928), .B2(new_n894), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n929), .A2(KEYINPUT118), .B1(new_n695), .B2(new_n452), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n926), .C1(new_n928), .C2(new_n894), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n906), .A2(new_n792), .A3(new_n793), .A4(new_n908), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n904), .B1(new_n933), .B2(new_n934), .ZN(G54));
  NAND4_X1  g749(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(new_n908), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n511), .ZN(new_n937));
  INV_X1    g751(.A(new_n904), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OR3_X1    g753(.A1(new_n936), .A2(KEYINPUT119), .A3(new_n511), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT119), .B1(new_n936), .B2(new_n511), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G60));
  INV_X1    g756(.A(new_n655), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n928), .B2(new_n894), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n938), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n901), .A2(new_n945), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n943), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND4_X1  g766(.A1(new_n882), .A2(new_n886), .A3(new_n680), .A4(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n882), .A2(new_n886), .A3(new_n952), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n938), .B(new_n953), .C1(new_n954), .C2(new_n384), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT61), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n524), .B2(new_n584), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n875), .B2(G953), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT121), .Z(new_n961));
  OAI21_X1  g775(.A(new_n910), .B1(G898), .B2(new_n344), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n250), .A2(new_n252), .ZN(new_n964));
  MUX2_X1   g778(.A(new_n507), .B(new_n351), .S(KEYINPUT19), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n690), .A2(new_n722), .A3(new_n747), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n771), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n765), .A2(new_n388), .A3(new_n742), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n970), .B(new_n769), .C1(new_n797), .C2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n798), .A2(new_n972), .A3(new_n806), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n968), .B1(new_n973), .B2(new_n344), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n766), .A2(new_n698), .A3(new_n699), .A4(new_n871), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n800), .A2(new_n975), .A3(new_n638), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  INV_X1    g791(.A(new_n969), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n717), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n704), .A2(new_n705), .ZN(new_n980));
  INV_X1    g794(.A(new_n716), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n701), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT62), .B(new_n969), .C1(new_n982), .C2(new_n712), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n976), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n786), .A2(new_n797), .ZN(new_n985));
  INV_X1    g799(.A(new_n806), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n344), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n974), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  AND2_X1   g806(.A1(G227), .A2(G900), .ZN(new_n993));
  OAI22_X1  g807(.A1(new_n974), .A2(new_n992), .B1(new_n344), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n988), .A2(KEYINPUT122), .A3(new_n966), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n991), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  NAND4_X1  g812(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n875), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT124), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n999), .A2(KEYINPUT125), .A3(new_n1002), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1005), .A2(new_n268), .A3(new_n247), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n973), .A2(new_n875), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n268), .A2(new_n247), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n904), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n270), .A2(new_n275), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1001), .B1(new_n1013), .B2(new_n707), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT126), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n900), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(G57));
endmodule


