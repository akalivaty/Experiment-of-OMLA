//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(G355));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G58), .C2(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n227), .B(new_n229), .C1(new_n219), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n223), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n206), .A2(new_n207), .ZN(new_n234));
  AOI22_X1  g0034(.A1(new_n231), .A2(KEYINPUT0), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n226), .B(new_n235), .C1(KEYINPUT0), .C2(new_n231), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  INV_X1    g0041(.A(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n214), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n213), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G226), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI211_X1 g0058(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT67), .B1(new_n268), .B2(G274), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n263), .A2(new_n270), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G238), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n265), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n265), .A2(new_n274), .A3(new_n281), .A4(new_n277), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n265), .A2(new_n277), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n281), .A4(new_n274), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(G169), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n279), .A2(G179), .A3(new_n282), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n283), .A2(new_n289), .A3(G169), .A4(new_n285), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n293), .A2(G77), .B1(new_n294), .B2(G50), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n223), .B2(G68), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n297), .A2(new_n232), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT11), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT69), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n222), .A2(G13), .A3(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  AND4_X1   g0104(.A1(new_n302), .A2(new_n303), .A3(new_n232), .A4(new_n297), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n222), .B2(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G68), .ZN(new_n308));
  INV_X1    g0108(.A(new_n303), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n202), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n301), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n291), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n312), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(G200), .A3(new_n285), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n279), .A2(G190), .A3(new_n282), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n292), .ZN(new_n319));
  NAND2_X1  g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G232), .A3(new_n255), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(G1698), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n323), .B2(new_n321), .C1(new_n324), .C2(new_n217), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n264), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n276), .A2(G244), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n274), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n307), .A2(G77), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT8), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G58), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT15), .B(G87), .Z(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n294), .B1(new_n293), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n223), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n299), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n332), .B(new_n342), .C1(G77), .C2(new_n303), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n331), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n313), .A2(new_n317), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n321), .A2(G222), .A3(new_n255), .ZN(new_n348));
  INV_X1    g0148(.A(G223), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n348), .B1(new_n340), .B2(new_n321), .C1(new_n324), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n264), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(new_n274), .C1(new_n242), .C2(new_n275), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(G179), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT68), .B1(new_n201), .B2(KEYINPUT8), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n333), .B2(G58), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n293), .B1(new_n208), .B2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n294), .A2(G150), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n299), .B1(new_n207), .B2(new_n309), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n299), .B1(new_n222), .B2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G50), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n352), .A2(new_n344), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n353), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n343), .B1(G200), .B2(new_n328), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n329), .A2(G190), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n361), .A2(new_n363), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(KEYINPUT9), .B1(G200), .B2(new_n352), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n352), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n371), .A2(new_n378), .A3(new_n373), .A4(new_n375), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n366), .B(new_n369), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  INV_X1    g0181(.A(new_n357), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n303), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n382), .B2(new_n362), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n203), .A2(new_n205), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n294), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n319), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n320), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT71), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n319), .A2(new_n223), .A3(new_n320), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n392), .A3(new_n391), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n298), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n401), .A3(new_n391), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(KEYINPUT72), .A3(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(G68), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n388), .A2(new_n389), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n385), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n269), .A2(new_n273), .B1(new_n275), .B2(new_n239), .ZN(new_n410));
  OAI211_X1 g0210(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT73), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT73), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n321), .A2(new_n413), .A3(G226), .A4(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n321), .A2(G223), .A3(new_n255), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n410), .B1(new_n417), .B2(new_n264), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n344), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n330), .B(new_n410), .C1(new_n417), .C2(new_n264), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n381), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n397), .A2(new_n392), .A3(new_n391), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n405), .B(KEYINPUT16), .C1(new_n423), .C2(new_n393), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n299), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT16), .B1(new_n404), .B2(new_n405), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n384), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n418), .A2(G179), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n344), .B2(new_n418), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT18), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(KEYINPUT74), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n429), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n381), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n418), .A2(G200), .ZN(new_n435));
  AOI211_X1 g0235(.A(G190), .B(new_n410), .C1(new_n417), .C2(new_n264), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT17), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n418), .A2(new_n372), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(G200), .B2(new_n418), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n409), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(new_n434), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT75), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n444), .A2(KEYINPUT75), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n347), .A2(new_n380), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n223), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n321), .A2(new_n223), .A3(G87), .A4(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n293), .A2(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n323), .A2(G20), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT88), .B1(new_n457), .B2(KEYINPUT23), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT88), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n323), .A4(G20), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n458), .A2(new_n461), .B1(KEYINPUT23), .B2(new_n457), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n455), .A2(new_n465), .A3(new_n456), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n299), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n222), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n298), .A2(new_n303), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n323), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT89), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n309), .B(new_n323), .C1(new_n473), .C2(KEYINPUT25), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(KEYINPUT25), .ZN(new_n475));
  XOR2_X1   g0275(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n468), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G294), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n264), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(G41), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n266), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n267), .A2(G1), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(G41), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G264), .A3(new_n263), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n486), .A2(new_n487), .ZN(new_n494));
  INV_X1    g0294(.A(new_n232), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n272), .B1(new_n495), .B2(new_n262), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n222), .A2(G45), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT78), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT78), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n500), .A3(new_n489), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n494), .A2(new_n496), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n344), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n330), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n478), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n471), .B1(new_n467), .B2(new_n299), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(G200), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .A4(new_n477), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n402), .A2(G107), .A3(new_n403), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT76), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n294), .A2(G77), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n323), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n514), .B(new_n515), .C1(new_n521), .C2(new_n223), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n223), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  INV_X1    g0323(.A(new_n515), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT76), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n513), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n299), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n303), .A2(G97), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n470), .A2(new_n218), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n321), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(G250), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n321), .A2(new_n540), .A3(G250), .A4(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n264), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n490), .A2(G257), .A3(new_n263), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n502), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(G190), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n527), .A2(new_n529), .A3(new_n531), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G200), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n544), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT80), .B1(new_n502), .B2(new_n544), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT81), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n528), .B(new_n530), .C1(new_n526), .C2(new_n299), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  INV_X1    g0356(.A(new_n551), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n544), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n543), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n555), .A2(new_n556), .A3(new_n560), .A4(new_n547), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n557), .A2(new_n543), .A3(new_n330), .A4(new_n558), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT82), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n552), .A2(new_n565), .A3(new_n330), .A4(new_n543), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n543), .A2(new_n546), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n344), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n562), .A2(new_n564), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n554), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n223), .B1(new_n260), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n518), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n223), .A2(G33), .A3(G97), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n574), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n321), .A2(new_n223), .A3(G68), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n298), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n470), .A2(new_n573), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n338), .A2(new_n303), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G238), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G116), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n264), .ZN(new_n586));
  AND2_X1   g0386(.A1(G33), .A2(G41), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n498), .B(G250), .C1(new_n587), .C2(new_n232), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n488), .A2(G274), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n586), .A2(G190), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n581), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n586), .A2(new_n592), .A3(new_n593), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n344), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n578), .A2(new_n580), .ZN(new_n601));
  INV_X1    g0401(.A(new_n338), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n470), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n588), .A2(KEYINPUT83), .A3(new_n589), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT83), .B1(new_n588), .B2(new_n589), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n330), .A3(new_n586), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n598), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n297), .A2(new_n232), .B1(G20), .B2(new_n213), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n536), .B(new_n223), .C1(G33), .C2(new_n218), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n612), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT20), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n611), .A2(KEYINPUT85), .A3(new_n612), .A4(KEYINPUT20), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n309), .A2(new_n213), .ZN(new_n621));
  OAI211_X1 g0421(.A(G116), .B(new_n469), .C1(new_n304), .C2(new_n305), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(G169), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n490), .A2(G270), .A3(new_n263), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n490), .A2(KEYINPUT84), .A3(G270), .A4(new_n263), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G303), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n324), .A2(new_n230), .B1(new_n631), .B2(new_n321), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n321), .A2(G257), .A3(new_n255), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n264), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n635), .A3(new_n502), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT21), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(KEYINPUT21), .A3(G169), .A4(new_n623), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT86), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(G169), .A3(new_n623), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n636), .A2(new_n330), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(new_n623), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n636), .A2(G200), .ZN(new_n645));
  INV_X1    g0445(.A(new_n623), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n645), .B(new_n646), .C1(new_n372), .C2(new_n636), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n610), .A2(new_n640), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n448), .A2(new_n512), .A3(new_n570), .A4(new_n648), .ZN(G372));
  NAND2_X1  g0449(.A1(new_n377), .A2(new_n379), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n443), .A2(new_n317), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n313), .B2(new_n346), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n422), .A2(new_n430), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n366), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n608), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n586), .A2(KEYINPUT90), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n585), .A2(new_n660), .A3(new_n264), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n604), .B2(new_n605), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n592), .A2(KEYINPUT91), .A3(new_n593), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n344), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(G200), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n658), .A2(new_n668), .B1(new_n669), .B2(new_n595), .ZN(new_n670));
  INV_X1    g0470(.A(new_n568), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n555), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n564), .A2(new_n566), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n670), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n569), .B2(new_n609), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n658), .A2(new_n668), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT92), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n507), .A2(new_n644), .A3(new_n640), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n554), .A2(new_n561), .A3(new_n569), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n511), .A2(new_n670), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n675), .A2(new_n676), .A3(new_n684), .A4(new_n677), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n657), .B1(new_n448), .B2(new_n687), .ZN(G369));
  AND2_X1   g0488(.A1(new_n640), .A2(new_n644), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n222), .A2(new_n223), .A3(G13), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT27), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT94), .B(G343), .Z(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT95), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n623), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n689), .A2(new_n647), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n689), .B2(new_n696), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT96), .ZN(new_n700));
  INV_X1    g0500(.A(new_n695), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n507), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n507), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n507), .A2(new_n511), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n478), .A2(new_n695), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n689), .A2(new_n695), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n704), .B2(new_n707), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n507), .A2(new_n695), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n714), .ZN(G399));
  NOR2_X1   g0515(.A1(new_n229), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n574), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n234), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n717), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n724));
  INV_X1    g0524(.A(new_n569), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT26), .A3(new_n670), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n674), .B1(new_n569), .B2(new_n609), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT98), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(KEYINPUT98), .B(new_n674), .C1(new_n569), .C2(new_n609), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT99), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n680), .A2(new_n681), .A3(new_n682), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n724), .A2(new_n731), .A3(new_n733), .A4(new_n677), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n723), .B1(new_n734), .B2(new_n701), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n686), .A2(new_n723), .A3(new_n701), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n630), .A2(new_n635), .A3(new_n502), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT97), .B1(new_n596), .B2(new_n492), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G179), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n493), .A2(new_n742), .A3(new_n606), .A4(new_n586), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n543), .A2(new_n546), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n738), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n596), .A2(new_n492), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n567), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(KEYINPUT30), .A3(new_n643), .A4(new_n740), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n552), .A2(new_n543), .B1(new_n662), .B2(new_n666), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n330), .A3(new_n503), .A4(new_n636), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n695), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n755), .A3(new_n695), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AND4_X1   g0557(.A1(new_n610), .A2(new_n640), .A3(new_n644), .A4(new_n647), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n705), .A3(new_n681), .A4(new_n701), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n737), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n735), .A2(new_n736), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n722), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n228), .A2(G20), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n717), .A2(G1), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n699), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n698), .ZN(new_n768));
  NAND2_X1  g0568(.A1(G20), .A2(G179), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT101), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n372), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n223), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(new_n372), .A3(new_n549), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n321), .B1(new_n777), .B2(G329), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n771), .A2(new_n330), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n778), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n372), .A2(new_n549), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n774), .B(new_n783), .C1(G326), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n770), .A2(new_n372), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G311), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n775), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G303), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n775), .A2(new_n372), .A3(G200), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT102), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n788), .A2(new_n549), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n796), .A2(G283), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n787), .A2(new_n790), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n218), .A2(new_n782), .B1(new_n785), .B2(new_n207), .ZN(new_n801));
  INV_X1    g0601(.A(new_n797), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n321), .B1(new_n802), .B2(new_n202), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G87), .C2(new_n792), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n777), .A2(G159), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  INV_X1    g0606(.A(new_n772), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G58), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n796), .A2(G107), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n789), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n340), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n800), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n232), .B1(G20), .B2(new_n344), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n250), .A2(G45), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n229), .A2(new_n321), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G45), .C2(new_n720), .ZN(new_n817));
  INV_X1    g0617(.A(new_n229), .ZN(new_n818));
  NAND3_X1  g0618(.A1(G355), .A2(new_n818), .A3(new_n321), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(G116), .C2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT100), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n814), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n813), .A2(new_n814), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n698), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n768), .B1(new_n765), .B2(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n346), .A2(new_n695), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n367), .A2(new_n368), .B1(new_n343), .B2(new_n695), .ZN(new_n832));
  INV_X1    g0632(.A(new_n346), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n687), .B2(new_n695), .ZN(new_n835));
  INV_X1    g0635(.A(new_n834), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n686), .A2(new_n701), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(new_n760), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n765), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n796), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n321), .B1(new_n776), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n781), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(new_n207), .C2(new_n791), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT103), .Z(new_n846));
  AOI22_X1  g0646(.A1(new_n797), .A2(G150), .B1(new_n786), .B2(G137), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  INV_X1    g0648(.A(G159), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n772), .C1(new_n849), .C2(new_n811), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT34), .Z(new_n851));
  NOR2_X1   g0651(.A1(new_n795), .A2(new_n573), .ZN(new_n852));
  INV_X1    g0652(.A(new_n321), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n791), .B2(new_n323), .ZN(new_n854));
  INV_X1    g0654(.A(G311), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n782), .A2(new_n218), .B1(new_n776), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G294), .C2(new_n807), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G116), .A2(new_n789), .B1(new_n797), .B2(G283), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n631), .C2(new_n785), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n846), .A2(new_n851), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n814), .A2(new_n821), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n860), .A2(new_n814), .B1(new_n340), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n862), .B(new_n766), .C1(new_n823), .C2(new_n836), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n840), .A2(new_n863), .ZN(G384));
  OAI21_X1  g0664(.A(new_n405), .B1(new_n423), .B2(new_n393), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n407), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n385), .B1(new_n400), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n692), .A2(G213), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n444), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n421), .A2(new_n867), .B1(new_n427), .B2(new_n437), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n409), .A2(new_n441), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT104), .C1(new_n421), .C2(new_n867), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(new_n868), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n427), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT37), .B1(new_n432), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n870), .B(KEYINPUT38), .C1(new_n877), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n875), .A2(new_n432), .A3(new_n880), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n881), .A2(new_n883), .B1(KEYINPUT37), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n653), .B2(new_n443), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n885), .A2(KEYINPUT106), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n872), .A2(new_n873), .ZN(new_n892));
  INV_X1    g0692(.A(new_n869), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n876), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n881), .A2(new_n883), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .A4(new_n870), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n757), .A2(new_n759), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n695), .A2(new_n312), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n313), .A2(new_n317), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n317), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n312), .B(new_n695), .C1(new_n291), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n836), .A4(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n870), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n894), .A2(KEYINPUT37), .B1(new_n881), .B2(new_n883), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n886), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n885), .ZN(new_n912));
  AOI221_X4 g0712(.A(new_n834), .B1(new_n903), .B2(new_n905), .C1(new_n757), .C2(new_n759), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n447), .A2(new_n901), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G330), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n447), .B1(new_n735), .B2(new_n736), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n657), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n313), .A2(new_n695), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT39), .B1(new_n891), .B2(new_n899), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n911), .B2(new_n885), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n906), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n837), .B2(new_n831), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n912), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n654), .A2(new_n868), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n921), .B(new_n931), .Z(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n222), .B2(new_n763), .ZN(new_n933));
  INV_X1    g0733(.A(new_n521), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n213), .B1(new_n934), .B2(KEYINPUT35), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n233), .C1(KEYINPUT35), .C2(new_n934), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n234), .A2(G77), .A3(new_n386), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(G50), .B2(new_n202), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n228), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n937), .A3(new_n940), .ZN(G367));
  NAND2_X1  g0741(.A1(new_n708), .A2(new_n710), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n681), .B1(new_n555), .B2(new_n701), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n725), .A2(new_n695), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT42), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n569), .B1(new_n943), .B2(new_n507), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n701), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n712), .A2(new_n950), .A3(new_n945), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT108), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n701), .A2(new_n581), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n670), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n677), .B2(new_n954), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT107), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n952), .A2(new_n953), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n953), .B1(new_n952), .B2(new_n958), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n952), .A2(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT108), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n952), .A2(new_n958), .A3(new_n953), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n709), .A2(new_n946), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n961), .A2(new_n966), .A3(KEYINPUT109), .A4(new_n967), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n967), .B1(new_n961), .B2(new_n966), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n764), .A2(G1), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n716), .B(KEYINPUT41), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT111), .B1(new_n714), .B2(new_n945), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT111), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n712), .A2(new_n946), .A3(new_n981), .A4(new_n713), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n979), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n713), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n942), .A2(new_n984), .A3(new_n945), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n981), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n714), .A2(KEYINPUT111), .A3(new_n945), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n978), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n714), .B2(new_n945), .ZN(new_n990));
  OAI211_X1 g0790(.A(KEYINPUT44), .B(new_n946), .C1(new_n712), .C2(new_n713), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n983), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n709), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n761), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n704), .A2(new_n711), .A3(new_n707), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(KEYINPUT113), .A3(new_n699), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n942), .B(KEYINPUT112), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n699), .A2(KEYINPUT113), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n699), .A2(KEYINPUT113), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n997), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n996), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n983), .A2(new_n988), .A3(new_n709), .A4(new_n992), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n995), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n977), .B1(new_n1008), .B2(new_n761), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n972), .B(new_n974), .C1(new_n975), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n321), .B1(new_n786), .B2(G311), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n631), .C2(new_n772), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT46), .B1(new_n792), .B2(G116), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n782), .A2(new_n323), .B1(new_n794), .B2(new_n218), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(G294), .C2(new_n797), .ZN(new_n1016));
  INV_X1    g0816(.A(G283), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1017), .B2(new_n811), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1013), .B(new_n1018), .C1(G317), .C2(new_n777), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT114), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n791), .A2(new_n201), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G50), .A2(new_n789), .B1(new_n797), .B2(G159), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n794), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G77), .A2(new_n1023), .B1(new_n781), .B2(G68), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G143), .A2(new_n786), .B1(new_n807), .B2(G150), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n853), .B1(new_n777), .B2(G137), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1020), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT47), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n765), .B1(new_n1029), .B2(new_n814), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n816), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n825), .B1(new_n818), .B2(new_n602), .C1(new_n246), .C2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n957), .A2(new_n827), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1010), .A2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n975), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n789), .A2(G303), .B1(new_n807), .B2(G317), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n855), .B2(new_n802), .C1(new_n773), .C2(new_n785), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT48), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n1017), .B2(new_n782), .C1(new_n779), .C2(new_n791), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n777), .A2(G326), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n321), .B1(new_n1023), .B2(G116), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n795), .A2(new_n218), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n207), .A2(new_n772), .B1(new_n785), .B2(new_n849), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G77), .B2(new_n792), .ZN(new_n1050));
  INV_X1    g0850(.A(G150), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n776), .A2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n853), .B(new_n1052), .C1(new_n338), .C2(new_n781), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G68), .A2(new_n789), .B1(new_n797), .B2(new_n357), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1047), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n718), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n818), .A3(new_n321), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n243), .A2(new_n267), .ZN(new_n1059));
  AOI211_X1 g0859(.A(G45), .B(new_n1057), .C1(G68), .C2(G77), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n336), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n336), .B2(G50), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n816), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1058), .B1(G107), .B2(new_n818), .C1(new_n1059), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1056), .A2(new_n814), .B1(new_n825), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n766), .C1(new_n708), .C2(new_n827), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n716), .B1(new_n1036), .B2(new_n761), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1037), .B(new_n1069), .C1(new_n1070), .C2(new_n1006), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n995), .A2(new_n1007), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1006), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n716), .A3(new_n1008), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n995), .A2(new_n975), .A3(new_n1007), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n945), .A2(new_n827), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n825), .B1(new_n218), .B2(new_n818), .C1(new_n253), .C2(new_n1031), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(KEYINPUT116), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G311), .A2(new_n807), .B1(new_n786), .B2(G317), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  AOI22_X1  g0883(.A1(G294), .A2(new_n789), .B1(new_n797), .B2(G303), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n853), .B1(new_n782), .B2(new_n213), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G322), .B2(new_n777), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n809), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n791), .A2(new_n1017), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n781), .A2(G77), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n811), .B2(new_n336), .C1(new_n207), .C2(new_n802), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n321), .B1(new_n791), .B2(new_n202), .C1(new_n848), .C2(new_n776), .ZN(new_n1091));
  OR3_X1    g0891(.A1(new_n1090), .A2(new_n852), .A3(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1051), .A2(new_n785), .B1(new_n772), .B2(new_n849), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n1087), .A2(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n765), .B1(new_n1095), .B2(new_n814), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1076), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1075), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT117), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1075), .A2(new_n1101), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(G390));
  AND3_X1   g0903(.A1(new_n760), .A2(new_n836), .A3(new_n906), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n837), .A2(new_n831), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n922), .B1(new_n1105), .B2(new_n906), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1106), .A2(new_n925), .A3(new_n923), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n832), .A2(new_n833), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n734), .A2(new_n701), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n927), .B1(new_n1110), .B2(new_n831), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1111), .A2(new_n922), .A3(new_n900), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1104), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n922), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n900), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1110), .A2(new_n831), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n1115), .C1(new_n1116), .C2(new_n927), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n923), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n925), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n928), .C2(new_n922), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n760), .A2(new_n836), .A3(new_n906), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n906), .B1(new_n760), .B2(new_n836), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1105), .B1(new_n1104), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n901), .A2(G330), .A3(new_n836), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n927), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1126), .A2(new_n1110), .A3(new_n1121), .A4(new_n831), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n447), .A2(G330), .A3(new_n901), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n919), .A2(new_n657), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n919), .A2(new_n657), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT118), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1113), .B(new_n1122), .C1(new_n1132), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1131), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(KEYINPUT118), .A3(new_n1134), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1107), .A2(new_n1112), .A3(new_n1104), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1121), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1141), .A3(new_n716), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1113), .A2(new_n975), .A3(new_n1122), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1113), .A2(new_n1122), .A3(KEYINPUT119), .A4(new_n975), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n853), .B1(new_n776), .B2(new_n779), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G87), .B2(new_n792), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n807), .A2(G116), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n786), .A2(G283), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1089), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n841), .B1(new_n323), .B2(new_n802), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(G97), .C2(new_n789), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT120), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G137), .A2(new_n797), .B1(new_n789), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n807), .A2(G132), .B1(G159), .B2(new_n781), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n785), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n853), .B1(new_n777), .B2(G125), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n207), .B2(new_n794), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT121), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n792), .A2(G150), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1160), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1154), .A2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(new_n814), .B1(new_n382), .B2(new_n861), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n766), .B(new_n1168), .C1(new_n1169), .C2(new_n823), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1142), .A2(new_n1147), .A3(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT122), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n908), .A2(new_n914), .A3(new_n737), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n931), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n891), .A4(new_n899), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n901), .A2(new_n836), .A3(new_n906), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n885), .B2(new_n911), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(G330), .C1(new_n1177), .C2(KEYINPUT40), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1178), .A2(new_n929), .A3(new_n926), .A4(new_n930), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n370), .A2(new_n868), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n650), .B2(new_n656), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n366), .B(new_n1180), .C1(new_n377), .C2(new_n379), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1182), .A2(new_n1183), .A3(KEYINPUT55), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT55), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1184), .A2(KEYINPUT56), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT56), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1174), .A2(new_n1179), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1172), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1188), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1174), .A2(new_n1179), .A3(new_n1188), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT122), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n1196), .A3(new_n975), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n861), .A2(new_n207), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n853), .B(new_n266), .C1(new_n340), .C2(new_n791), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n794), .A2(new_n201), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G283), .B2(new_n777), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n202), .B2(new_n782), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1199), .B(new_n1202), .C1(G107), .C2(new_n807), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G97), .A2(new_n797), .B1(new_n789), .B2(new_n338), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n213), .C2(new_n785), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G132), .A2(new_n797), .B1(new_n789), .B2(G137), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n807), .A2(G128), .B1(G150), .B2(new_n781), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1156), .A2(new_n792), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n786), .A2(G125), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1210), .A2(KEYINPUT59), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT59), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G33), .B1(new_n1023), .B2(G159), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G41), .B1(new_n777), .B2(G124), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n207), .B1(new_n256), .B2(G41), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1206), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n765), .B1(new_n1218), .B2(new_n814), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1198), .B(new_n1219), .C1(new_n1193), .C2(new_n823), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1197), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1136), .A2(new_n1133), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n1191), .A3(new_n1196), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1136), .A2(new_n1133), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n717), .B1(new_n1226), .B2(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1221), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(G375));
  OAI22_X1  g1029(.A1(new_n782), .A2(new_n207), .B1(new_n776), .B2(new_n1159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n853), .B(new_n1230), .C1(G159), .C2(new_n792), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n797), .A2(new_n1156), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n789), .A2(G150), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n785), .A2(new_n842), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1200), .B(new_n1234), .C1(G137), .C2(new_n807), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n853), .B1(new_n791), .B2(new_n218), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n782), .A2(new_n602), .B1(new_n631), .B2(new_n776), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(G294), .C2(new_n786), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n796), .A2(G77), .B1(G116), .B2(new_n797), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n1017), .C2(new_n772), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n811), .A2(new_n323), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1236), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT123), .Z(new_n1244));
  AOI21_X1  g1044(.A(new_n765), .B1(new_n1244), .B2(new_n814), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n821), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n906), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n202), .B2(new_n861), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1134), .B2(new_n975), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1137), .A2(new_n1138), .A3(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(new_n977), .ZN(G381));
  NAND4_X1  g1052(.A1(new_n1010), .A2(new_n1034), .A3(new_n1102), .A4(new_n1100), .ZN(new_n1253));
  OR3_X1    g1053(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1254));
  OR3_X1    g1054(.A1(new_n1253), .A2(G381), .A3(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(KEYINPUT124), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1170), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1142), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G375), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1256), .A2(new_n1257), .A3(new_n1265), .ZN(G407));
  INV_X1    g1066(.A(new_n693), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(G213), .ZN(new_n1268));
  XOR2_X1   g1068(.A(new_n1268), .B(KEYINPUT126), .Z(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  NAND2_X1  g1071(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1221), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(G378), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n975), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1220), .B(new_n1275), .C1(new_n1223), .C2(new_n977), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1262), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1261), .B1(new_n1260), .B2(new_n1142), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1274), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1269), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1251), .A2(KEYINPUT60), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n717), .B1(new_n1250), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1282), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1249), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1282), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT127), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G384), .B(new_n1249), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1280), .A2(new_n1281), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1249), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n840), .A3(new_n863), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1269), .A2(G2897), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1293), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1301), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1228), .A2(G378), .B1(new_n1263), .B2(new_n1276), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1302), .B(new_n1304), .C1(new_n1305), .C2(new_n1269), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1269), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1295), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1297), .A2(new_n1298), .A3(new_n1306), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1008), .A2(new_n761), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n975), .B1(new_n1311), .B2(new_n976), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n970), .A2(new_n971), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n973), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1034), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1075), .A2(new_n1101), .A3(new_n1098), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1101), .B1(new_n1075), .B2(new_n1098), .ZN(new_n1317));
  OAI22_X1  g1117(.A1(new_n1314), .A2(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(G393), .B(G396), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1253), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1253), .B2(new_n1318), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1310), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1304), .A2(new_n1302), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT63), .B1(new_n1325), .B2(new_n1307), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1296), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1281), .A4(new_n1295), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1322), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1327), .A2(new_n1329), .A3(new_n1298), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1330), .ZN(G405));
  NOR2_X1   g1131(.A1(new_n1264), .A2(new_n1228), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1274), .ZN(new_n1333));
  OR3_X1    g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1295), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1295), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1323), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1334), .A2(new_n1322), .A3(new_n1335), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


