//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(new_n461), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g054(.A1(new_n463), .A2(new_n465), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n463), .A2(new_n465), .A3(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT70), .ZN(G162));
  NAND3_X1  g063(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n461), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n461), .A2(G102), .A3(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT71), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  INV_X1    g070(.A(new_n490), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n471), .B2(G126), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n495), .B(new_n492), .C1(new_n497), .C2(new_n461), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT72), .A4(new_n461), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n483), .A2(KEYINPUT72), .A3(KEYINPUT4), .A4(G138), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n494), .A2(new_n498), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT75), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI211_X1 g084(.A(G50), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n512), .B(new_n514), .C1(new_n508), .C2(new_n509), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n507), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(G88), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n507), .B1(new_n521), .B2(new_n510), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n512), .A2(new_n514), .A3(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n512), .A2(new_n514), .A3(new_n527), .A4(G62), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n506), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(new_n510), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n517), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(KEYINPUT75), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n531), .A2(new_n536), .ZN(G166));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT76), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(G63), .A2(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n508), .A2(new_n509), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(new_n519), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n511), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G51), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n541), .A2(new_n549), .ZN(G168));
  AOI22_X1  g125(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  INV_X1    g130(.A(G90), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n554), .A2(new_n555), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(G171));
  AOI22_X1  g133(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n552), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  INV_X1    g136(.A(G81), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n554), .A2(new_n561), .B1(new_n515), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(KEYINPUT77), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n560), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  AOI22_X1  g150(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n576), .A2(new_n552), .B1(new_n577), .B2(new_n515), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n547), .A2(KEYINPUT9), .A3(G53), .ZN(new_n579));
  AOI21_X1  g154(.A(KEYINPUT9), .B1(new_n547), .B2(G53), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  OR2_X1    g158(.A1(new_n539), .A2(new_n540), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n539), .A2(new_n540), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n584), .A2(new_n548), .A3(new_n546), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G286));
  INV_X1    g166(.A(G166), .ZN(G303));
  OAI21_X1  g167(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n520), .A2(G49), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n515), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(G288));
  NAND3_X1  g173(.A1(new_n519), .A2(new_n520), .A3(G86), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n520), .A2(G48), .A3(G543), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n552), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n552), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT81), .Z(new_n607));
  INV_X1    g182(.A(new_n515), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT82), .B(G85), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n547), .A2(G47), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n515), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n519), .A2(G66), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(new_n547), .B2(G54), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT84), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n615), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(new_n626), .A3(new_n621), .ZN(new_n627));
  AND2_X1   g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n613), .B1(new_n628), .B2(G868), .ZN(G284));
  OAI21_X1  g204(.A(new_n613), .B1(new_n628), .B2(G868), .ZN(G321));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(G299), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n590), .B2(new_n631), .ZN(G297));
  OAI21_X1  g208(.A(new_n632), .B1(new_n590), .B2(new_n631), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n628), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n481), .A2(G123), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n483), .A2(G135), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n648));
  NOR3_X1   g223(.A1(new_n464), .A2(new_n462), .A3(G2105), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(KEYINPUT86), .A2(G2100), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT13), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(G14), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n676), .A3(KEYINPUT17), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT19), .Z(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n689), .A2(new_n690), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n690), .C2(new_n689), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G1981), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  OR2_X1    g276(.A1(G29), .A2(G32), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G129), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT98), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n483), .A2(G141), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n703), .A2(new_n705), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n702), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1996), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(G1996), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n711), .A2(G27), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n504), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G2078), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(G171), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G5), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n719), .A2(new_n723), .A3(new_n724), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(G160), .A2(G29), .ZN(new_n730));
  AND2_X1   g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  NOR2_X1   g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n711), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(G2084), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n483), .A2(G139), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI22_X1  g313(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT97), .Z(new_n740));
  OAI211_X1 g315(.A(new_n736), .B(new_n738), .C1(new_n740), .C2(new_n461), .ZN(new_n741));
  MUX2_X1   g316(.A(G33), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  OR2_X1    g318(.A1(G16), .A2(G21), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n586), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT30), .B(G28), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n746), .A2(new_n747), .B1(new_n711), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n645), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  OAI211_X1 g327(.A(G1966), .B(new_n744), .C1(new_n586), .C2(new_n745), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n749), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n726), .A2(new_n727), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n755), .B1(new_n754), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n730), .A2(G2084), .A3(new_n733), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n735), .A2(new_n743), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n762));
  INV_X1    g337(.A(new_n760), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n729), .A2(new_n763), .A3(new_n734), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n764), .A2(new_n765), .A3(new_n743), .A4(new_n759), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n711), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n711), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(G2090), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n745), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n569), .B2(new_n745), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1341), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n771), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n762), .A2(new_n766), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n481), .A2(G119), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n483), .A2(G131), .ZN(new_n779));
  NOR2_X1   g354(.A1(G95), .A2(G2105), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G25), .B(new_n782), .S(G29), .Z(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT35), .B(G1991), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT90), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G290), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n745), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n745), .B2(G24), .ZN(new_n789));
  INV_X1    g364(.A(G1986), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n745), .A2(G6), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G305), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT32), .B(G1981), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n745), .A2(G23), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n596), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n608), .A2(G87), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n801), .A2(KEYINPUT92), .A3(new_n594), .A4(new_n593), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n803), .B2(new_n745), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT33), .B(G1976), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT93), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n745), .B1(new_n531), .B2(new_n536), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(G1971), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n808), .A2(G1971), .A3(new_n809), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n797), .B(new_n807), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  INV_X1    g391(.A(new_n812), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n810), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n818), .A2(KEYINPUT94), .A3(new_n807), .A4(new_n797), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n815), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n792), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n792), .B1(new_n823), .B2(new_n824), .C1(new_n820), .C2(new_n821), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n777), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n745), .A2(G20), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G299), .B2(G16), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1956), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n711), .A2(G26), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n481), .A2(G128), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n483), .A2(G140), .ZN(new_n836));
  NOR2_X1   g411(.A1(G104), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n834), .B1(new_n839), .B2(G29), .ZN(new_n840));
  MUX2_X1   g415(.A(new_n834), .B(new_n840), .S(KEYINPUT28), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G2067), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n745), .A2(G4), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n628), .B2(new_n745), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT96), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G1348), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n828), .A2(new_n833), .A3(new_n842), .A4(new_n847), .ZN(G150));
  NAND2_X1  g423(.A1(G150), .A2(KEYINPUT102), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n846), .B(new_n777), .C1(new_n826), .C2(new_n827), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n833), .A4(new_n842), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(G311));
  AOI22_X1  g428(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n552), .ZN(new_n855));
  INV_X1    g430(.A(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n554), .A2(new_n856), .B1(new_n515), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n568), .B(new_n859), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n628), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n635), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n865), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n862), .B1(new_n868), .B2(G860), .ZN(G145));
  XNOR2_X1  g444(.A(new_n782), .B(new_n710), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n478), .B(KEYINPUT69), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n645), .ZN(new_n872));
  NAND2_X1  g447(.A1(G160), .A2(new_n750), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(G162), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G162), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n489), .A2(new_n490), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G2105), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n503), .A2(new_n879), .A3(new_n502), .A4(new_n492), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n650), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G162), .ZN(new_n883));
  INV_X1    g458(.A(new_n873), .ZN(new_n884));
  NOR2_X1   g459(.A1(G160), .A2(new_n750), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n870), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n874), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n877), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n882), .B1(new_n877), .B2(new_n888), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n741), .B(new_n839), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n481), .A2(G130), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n483), .A2(G142), .ZN(new_n893));
  NOR2_X1   g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n891), .B(new_n896), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n889), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n898), .A2(new_n899), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(G395));
  NAND2_X1  g482(.A1(G303), .A2(new_n803), .ZN(new_n908));
  NAND3_X1  g483(.A1(G166), .A2(new_n800), .A3(new_n802), .ZN(new_n909));
  AOI21_X1  g484(.A(G305), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(G305), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n787), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n914), .A2(new_n910), .A3(G290), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n863), .B(new_n637), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n625), .A2(new_n621), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n581), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n921), .B2(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n927), .B(new_n928), .C1(new_n913), .C2(new_n915), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n918), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n926), .B1(new_n918), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n860), .A2(new_n631), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  XNOR2_X1  g510(.A(G295), .B(new_n935), .ZN(G331));
  OAI21_X1  g511(.A(G171), .B1(new_n588), .B2(new_n589), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n937), .A2(KEYINPUT106), .B1(new_n586), .B2(G171), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT78), .ZN(new_n939));
  NAND2_X1  g514(.A1(G168), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G301), .B1(new_n940), .B2(new_n587), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n863), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n921), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n568), .B(new_n860), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n941), .A2(new_n942), .B1(G168), .B2(G301), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n937), .A2(KEYINPUT106), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n944), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n944), .A2(new_n949), .B1(new_n922), .B2(new_n923), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n916), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n944), .A2(new_n949), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n924), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n921), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g532(.A(G290), .B1(new_n914), .B2(new_n910), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n911), .A2(new_n787), .A3(new_n912), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n953), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n961), .A3(new_n900), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n915), .B2(new_n913), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n952), .A2(new_n916), .ZN(new_n966));
  AND4_X1   g541(.A1(KEYINPUT43), .A2(new_n965), .A3(new_n900), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT108), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(new_n963), .A3(new_n900), .A4(new_n966), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(new_n972), .A3(KEYINPUT43), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n478), .A2(G40), .A3(new_n976), .A4(new_n880), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G2067), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n494), .A2(new_n498), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n503), .A2(new_n502), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n983), .B(new_n468), .C1(new_n473), .C2(new_n477), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n880), .A2(new_n985), .A3(new_n976), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1348), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n866), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n978), .B(new_n628), .C1(new_n988), .C2(new_n989), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT60), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT61), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n504), .B2(new_n976), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n492), .B1(new_n497), .B2(new_n461), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n976), .C1(new_n980), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n984), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT56), .B(G2072), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n504), .A2(new_n985), .A3(new_n976), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n976), .B1(new_n980), .B2(new_n996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n984), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1956), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n999), .A2(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n581), .B(KEYINPUT57), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n994), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n984), .A2(new_n997), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n981), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1012), .A3(new_n1000), .ZN(new_n1013));
  AND4_X1   g588(.A1(new_n994), .A2(new_n1009), .A3(new_n1007), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(new_n1012), .A3(new_n716), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT58), .B(G1341), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n977), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT59), .B1(new_n1019), .B2(new_n569), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(new_n568), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n990), .A2(new_n1024), .A3(new_n628), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n993), .A2(new_n1015), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1006), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1007), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n991), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n995), .A2(new_n998), .A3(G2078), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n985), .B1(new_n504), .B2(new_n976), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n478), .A2(G40), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n986), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1032), .A2(KEYINPUT53), .B1(new_n1035), .B2(G1961), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n984), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n997), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n984), .A2(new_n1037), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2078), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1042), .B2(G2078), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NOR4_X1   g621(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G171), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n999), .A2(new_n722), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1039), .B(new_n984), .C1(new_n981), .C2(new_n1011), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n722), .A2(KEYINPUT53), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n988), .A2(new_n727), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1050), .A2(new_n1054), .A3(G301), .A4(new_n1055), .ZN(new_n1056));
  AND4_X1   g631(.A1(KEYINPUT123), .A2(new_n1048), .A3(KEYINPUT54), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(KEYINPUT112), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n531), .A2(new_n536), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(KEYINPUT112), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1061), .B(new_n1063), .Z(new_n1064));
  INV_X1    g639(.A(G1971), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n995), .B2(new_n998), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT111), .B(G2090), .Z(new_n1068));
  NAND4_X1  g643(.A1(new_n1001), .A2(new_n984), .A3(new_n1003), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1064), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n519), .A2(G61), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G73), .A2(G543), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n552), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n599), .A2(new_n600), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1981), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT116), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n602), .A2(new_n1083), .A3(G1981), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1074), .B(new_n1075), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(KEYINPUT116), .A3(new_n1081), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1083), .B1(new_n602), .B2(G1981), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1088), .A2(new_n1089), .B1(G1981), .B2(new_n602), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT49), .B1(new_n1090), .B2(KEYINPUT117), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1002), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1058), .B1(new_n1092), .B2(new_n984), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n803), .A2(G1976), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n803), .A2(KEYINPUT115), .A3(G1976), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1093), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT52), .ZN(new_n1100));
  INV_X1    g675(.A(G1976), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT52), .B1(G288), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(new_n1097), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1094), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n982), .A2(new_n987), .A3(new_n984), .A4(new_n1068), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1058), .B1(new_n1105), .B2(new_n1066), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1061), .B(new_n1063), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1073), .B(new_n1104), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1057), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1048), .A2(KEYINPUT54), .A3(new_n1056), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1051), .A2(new_n747), .ZN(new_n1116));
  INV_X1    g691(.A(G2084), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n982), .A2(new_n987), .A3(new_n1117), .A4(new_n984), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(G8), .A3(new_n586), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n586), .A2(G8), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1035), .A2(new_n1117), .B1(new_n1051), .B2(new_n747), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1123), .B(new_n1124), .C1(new_n1125), .C2(new_n1058), .ZN(new_n1126));
  OAI211_X1 g701(.A(G8), .B(new_n1122), .C1(new_n1119), .C2(new_n586), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1038), .A2(new_n1039), .A3(new_n997), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1041), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1043), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1045), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1050), .A2(new_n1133), .A3(G301), .A4(new_n1055), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1036), .A2(new_n1053), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(G301), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1120), .A2(new_n1129), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1031), .A2(new_n1112), .A3(new_n1115), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1129), .A2(new_n1120), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT62), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1111), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1135), .A2(G301), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1129), .A2(new_n1144), .A3(new_n1120), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1094), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1125), .A2(new_n1058), .A3(G286), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1073), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT114), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1148), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1093), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1158));
  INV_X1    g733(.A(G288), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(new_n1101), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1085), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1119), .A2(G8), .A3(new_n590), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1164), .A2(new_n1148), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1163), .B1(new_n1166), .B2(new_n1149), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1147), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(new_n1104), .A3(new_n1150), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1162), .B1(new_n1170), .B2(KEYINPUT63), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT118), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(G8), .A3(new_n1070), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n1174), .B2(new_n1064), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1175), .A2(new_n1150), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT119), .B(new_n1171), .C1(new_n1176), .C2(new_n1148), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1139), .A2(new_n1146), .A3(new_n1168), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1179), .A2(KEYINPUT109), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(KEYINPUT109), .ZN(new_n1181));
  OAI211_X1 g756(.A(G1996), .B(new_n710), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT110), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1179), .A2(new_n716), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n710), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1179), .B(KEYINPUT109), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n839), .B(G2067), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1187), .A2(KEYINPUT110), .A3(G1996), .A4(new_n710), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n782), .A2(new_n784), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n782), .A2(new_n784), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1187), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1184), .A2(new_n1189), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G290), .B(G1986), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1179), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1178), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1194), .A2(KEYINPUT125), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1194), .A2(KEYINPUT125), .ZN(new_n1200));
  NOR4_X1   g775(.A1(G290), .A2(G1986), .A3(new_n1039), .A4(new_n1034), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1191), .B(KEYINPUT124), .ZN(new_n1204));
  AND4_X1   g779(.A1(new_n1189), .A2(new_n1184), .A3(new_n1190), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n839), .A2(G2067), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1187), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1187), .B1(new_n710), .B2(new_n1188), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1185), .B(KEYINPUT46), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT47), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1207), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(KEYINPUT126), .B1(new_n1203), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1200), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1202), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1214), .A2(new_n1215), .A3(new_n1198), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1216), .A2(new_n1217), .A3(new_n1211), .A4(new_n1207), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1213), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1197), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1197), .A2(KEYINPUT127), .A3(new_n1219), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g799(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n1226));
  NOR2_X1   g800(.A1(G401), .A2(G227), .ZN(new_n1227));
  AND2_X1   g801(.A1(new_n901), .A2(new_n1227), .ZN(new_n1228));
  AND4_X1   g802(.A1(G319), .A2(new_n1226), .A3(new_n700), .A4(new_n1228), .ZN(G308));
  NAND4_X1  g803(.A1(new_n1226), .A2(G319), .A3(new_n700), .A4(new_n1228), .ZN(G225));
endmodule


