

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(n364), .B(KEYINPUT45), .ZN(n365) );
  XOR2_X1 U323 ( .A(n553), .B(KEYINPUT36), .Z(n583) );
  INV_X1 U324 ( .A(G190GAT), .ZN(n453) );
  XNOR2_X1 U325 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U326 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n291) );
  XNOR2_X1 U328 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n290) );
  XNOR2_X1 U329 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U330 ( .A(KEYINPUT17), .B(n292), .Z(n407) );
  XOR2_X1 U331 ( .A(G176GAT), .B(KEYINPUT86), .Z(n294) );
  XNOR2_X1 U332 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n305) );
  XOR2_X1 U334 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n296) );
  XOR2_X1 U335 ( .A(G190GAT), .B(G134GAT), .Z(n353) );
  XOR2_X1 U336 ( .A(G120GAT), .B(G71GAT), .Z(n311) );
  XNOR2_X1 U337 ( .A(n353), .B(n311), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U339 ( .A(n297), .B(G99GAT), .Z(n303) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n298), .B(G127GAT), .ZN(n434) );
  XOR2_X1 U342 ( .A(n434), .B(G169GAT), .Z(n300) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U347 ( .A(n305), .B(n304), .Z(n306) );
  XOR2_X1 U348 ( .A(n407), .B(n306), .Z(n460) );
  XNOR2_X1 U349 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n414) );
  XOR2_X1 U350 ( .A(G92GAT), .B(G64GAT), .Z(n308) );
  XNOR2_X1 U351 ( .A(G176GAT), .B(KEYINPUT76), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(G204GAT), .B(n309), .Z(n408) );
  XOR2_X1 U354 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n313) );
  XNOR2_X1 U355 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n310), .B(KEYINPUT71), .ZN(n339) );
  XNOR2_X1 U357 ( .A(n311), .B(n339), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n408), .B(n314), .ZN(n324) );
  XOR2_X1 U360 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n316) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n317), .B(KEYINPUT72), .Z(n322) );
  XOR2_X1 U364 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n421) );
  XNOR2_X1 U367 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n320), .B(KEYINPUT74), .ZN(n352) );
  XNOR2_X1 U369 ( .A(n421), .B(n352), .ZN(n321) );
  XNOR2_X1 U370 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U371 ( .A(n324), .B(n323), .Z(n457) );
  INV_X1 U372 ( .A(n457), .ZN(n574) );
  XOR2_X1 U373 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n326) );
  XNOR2_X1 U374 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n338) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G71GAT), .Z(n328) );
  XNOR2_X1 U377 ( .A(G183GAT), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n336) );
  XOR2_X1 U379 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n330) );
  XNOR2_X1 U380 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U382 ( .A(G64GAT), .B(G155GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(G22GAT), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n334), .B(n333), .Z(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .Z(n369) );
  XOR2_X1 U389 ( .A(n339), .B(n369), .Z(n341) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U392 ( .A(n343), .B(n342), .Z(n579) );
  INV_X1 U393 ( .A(n579), .ZN(n486) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n345) );
  XNOR2_X1 U395 ( .A(G50GAT), .B(KEYINPUT65), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n363) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(G92GAT), .Z(n347) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G218GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n349) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(G162GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U403 ( .A(n351), .B(n350), .Z(n361) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n355) );
  AND2_X1 U405 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n357) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G29GAT), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U410 ( .A(KEYINPUT7), .B(n358), .Z(n380) );
  XNOR2_X1 U411 ( .A(n359), .B(n380), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X2 U413 ( .A(n363), .B(n362), .ZN(n553) );
  NOR2_X1 U414 ( .A1(n486), .A2(n583), .ZN(n364) );
  INV_X1 U415 ( .A(n365), .ZN(n366) );
  NOR2_X1 U416 ( .A1(n574), .A2(n366), .ZN(n367) );
  XNOR2_X1 U417 ( .A(n367), .B(KEYINPUT113), .ZN(n383) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G36GAT), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n368), .B(G8GAT), .ZN(n402) );
  XOR2_X1 U420 ( .A(n369), .B(n402), .Z(n371) );
  XNOR2_X1 U421 ( .A(G113GAT), .B(G197GAT), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n376) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(G22GAT), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n372), .B(G141GAT), .ZN(n422) );
  XOR2_X1 U425 ( .A(n422), .B(KEYINPUT66), .Z(n374) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U428 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U429 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n378) );
  XNOR2_X1 U430 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U433 ( .A(n382), .B(n381), .Z(n500) );
  XOR2_X1 U434 ( .A(n500), .B(KEYINPUT70), .Z(n557) );
  NOR2_X1 U435 ( .A1(n383), .A2(n557), .ZN(n385) );
  INV_X1 U436 ( .A(KEYINPUT114), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n393) );
  INV_X1 U438 ( .A(n500), .ZN(n571) );
  XNOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n386) );
  XOR2_X1 U440 ( .A(n386), .B(n574), .Z(n548) );
  NAND2_X1 U441 ( .A1(n571), .A2(n548), .ZN(n388) );
  XNOR2_X1 U442 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  NAND2_X1 U444 ( .A1(n389), .A2(n486), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n553), .A2(n390), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT47), .B(n391), .ZN(n392) );
  NAND2_X1 U447 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U448 ( .A(KEYINPUT48), .B(n394), .ZN(n528) );
  XOR2_X1 U449 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n396) );
  XNOR2_X1 U450 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U452 ( .A(n397), .B(KEYINPUT90), .Z(n399) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(G211GAT), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n428) );
  XOR2_X1 U455 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n401) );
  XNOR2_X1 U456 ( .A(G190GAT), .B(KEYINPUT93), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT95), .B(n402), .Z(n404) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U461 ( .A(n406), .B(n405), .Z(n411) );
  INV_X1 U462 ( .A(n407), .ZN(n409) );
  XOR2_X1 U463 ( .A(n409), .B(n408), .Z(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U465 ( .A(n428), .B(n412), .Z(n518) );
  AND2_X1 U466 ( .A1(n528), .A2(n518), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n415) );
  INV_X1 U468 ( .A(n415), .ZN(n568) );
  XOR2_X1 U469 ( .A(G204GAT), .B(KEYINPUT22), .Z(n417) );
  NAND2_X1 U470 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n420) );
  XOR2_X1 U472 ( .A(G155GAT), .B(KEYINPUT2), .Z(n419) );
  XNOR2_X1 U473 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n437) );
  XOR2_X1 U475 ( .A(n420), .B(n437), .Z(n424) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n426) );
  XNOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U481 ( .A(n428), .B(n427), .Z(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n464) );
  XOR2_X1 U483 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n436) );
  XOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n432) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G57GAT), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n441) );
  XOR2_X1 U489 ( .A(n437), .B(G134GAT), .Z(n439) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U492 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U493 ( .A(G85GAT), .B(G148GAT), .Z(n443) );
  XNOR2_X1 U494 ( .A(G141GAT), .B(G120GAT), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n527) );
  INV_X1 U498 ( .A(n527), .ZN(n567) );
  AND2_X1 U499 ( .A1(n464), .A2(n567), .ZN(n447) );
  NAND2_X1 U500 ( .A1(n568), .A2(n447), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  NOR2_X1 U503 ( .A1(n460), .A2(n450), .ZN(n452) );
  INV_X1 U504 ( .A(KEYINPUT123), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n563) );
  NAND2_X1 U506 ( .A1(n563), .A2(n553), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n477) );
  NAND2_X1 U509 ( .A1(n557), .A2(n457), .ZN(n489) );
  XOR2_X1 U510 ( .A(n518), .B(KEYINPUT97), .Z(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n458), .Z(n467) );
  XOR2_X1 U512 ( .A(KEYINPUT28), .B(n464), .Z(n522) );
  NOR2_X1 U513 ( .A1(n467), .A2(n522), .ZN(n530) );
  NAND2_X1 U514 ( .A1(n460), .A2(n530), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n459), .A2(n527), .ZN(n471) );
  INV_X1 U516 ( .A(n460), .ZN(n529) );
  NAND2_X1 U517 ( .A1(n518), .A2(n529), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n464), .A2(n461), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n527), .A2(n463), .ZN(n469) );
  NOR2_X1 U521 ( .A1(n529), .A2(n464), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n569) );
  INV_X1 U524 ( .A(n467), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n569), .A2(n468), .ZN(n542) );
  NAND2_X1 U526 ( .A1(n469), .A2(n542), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n485) );
  INV_X1 U528 ( .A(n485), .ZN(n475) );
  OR2_X1 U529 ( .A1(n486), .A2(n553), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT83), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT16), .B(n473), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n502) );
  NOR2_X1 U533 ( .A1(n489), .A2(n502), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n483), .A2(n527), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n483), .A2(n518), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U540 ( .A1(n483), .A2(n529), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n522), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U545 ( .A1(n583), .A2(n485), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT37), .B(n488), .Z(n515) );
  NOR2_X1 U548 ( .A1(n515), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n490), .ZN(n498) );
  NAND2_X1 U550 ( .A1(n498), .A2(n527), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n498), .A2(n518), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n496) );
  NAND2_X1 U557 ( .A1(n498), .A2(n529), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n497), .Z(G1330GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n522), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n504) );
  XNOR2_X1 U563 ( .A(KEYINPUT104), .B(n548), .ZN(n559) );
  NAND2_X1 U564 ( .A1(n500), .A2(n559), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT105), .B(n501), .Z(n514) );
  NOR2_X1 U566 ( .A1(n514), .A2(n502), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n511), .A2(n527), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U571 ( .A1(n511), .A2(n518), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n529), .A2(n511), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n522), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(n516), .Z(n523) );
  NAND2_X1 U582 ( .A1(n527), .A2(n523), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT110), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U595 ( .A1(n541), .A2(n531), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n538), .A2(n557), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U599 ( .A1(n538), .A2(n559), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n579), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n553), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT116), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n571), .A2(n554), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(KEYINPUT52), .B(n547), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U619 ( .A1(n579), .A2(n554), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U627 ( .A1(n559), .A2(n563), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n579), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n573) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n582) );
  INV_X1 U637 ( .A(n582), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n580), .A2(n571), .ZN(n572) );
  XOR2_X1 U639 ( .A(n573), .B(n572), .Z(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U641 ( .A1(n580), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

