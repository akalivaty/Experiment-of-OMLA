

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745;

  NOR2_X1 U372 ( .A1(n708), .A2(n717), .ZN(n366) );
  NOR2_X1 U373 ( .A1(n659), .A2(n657), .ZN(n583) );
  OR2_X1 U374 ( .A1(n714), .A2(G902), .ZN(n399) );
  INV_X1 U375 ( .A(G953), .ZN(n731) );
  NOR2_X1 U376 ( .A1(n628), .A2(n717), .ZN(n631) );
  XNOR2_X2 U377 ( .A(n418), .B(G119), .ZN(n456) );
  XNOR2_X2 U378 ( .A(n491), .B(n414), .ZN(n445) );
  XNOR2_X2 U379 ( .A(n416), .B(G143), .ZN(n491) );
  XOR2_X2 U380 ( .A(G122), .B(G104), .Z(n505) );
  XNOR2_X2 U381 ( .A(n568), .B(n455), .ZN(n670) );
  XNOR2_X2 U382 ( .A(n454), .B(G469), .ZN(n568) );
  XNOR2_X2 U383 ( .A(n399), .B(n470), .ZN(n666) );
  NOR2_X1 U384 ( .A1(n618), .A2(n419), .ZN(n359) );
  NOR2_X1 U385 ( .A1(n643), .A2(n574), .ZN(n575) );
  INV_X1 U386 ( .A(n691), .ZN(n679) );
  INV_X1 U387 ( .A(G110), .ZN(n418) );
  INV_X1 U388 ( .A(G128), .ZN(n416) );
  AND2_X2 U389 ( .A1(n400), .A2(n372), .ZN(n710) );
  NAND2_X1 U390 ( .A1(n375), .A2(n371), .ZN(n400) );
  XNOR2_X1 U391 ( .A(n614), .B(n405), .ZN(n653) );
  XNOR2_X1 U392 ( .A(n526), .B(n525), .ZN(n585) );
  NOR2_X1 U393 ( .A1(G902), .A2(n698), .ZN(n454) );
  XNOR2_X1 U394 ( .A(n370), .B(G146), .ZN(n460) );
  XNOR2_X1 U395 ( .A(n415), .B(KEYINPUT65), .ZN(n414) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n514) );
  OR2_X1 U397 ( .A1(G902), .A2(G237), .ZN(n476) );
  XNOR2_X1 U398 ( .A(n487), .B(KEYINPUT21), .ZN(n562) );
  NAND2_X1 U399 ( .A1(n616), .A2(n651), .ZN(n617) );
  INV_X1 U400 ( .A(n652), .ZN(n616) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n609) );
  AND2_X1 U402 ( .A1(n608), .A2(n357), .ZN(n361) );
  AND2_X1 U403 ( .A1(n394), .A2(n564), .ZN(n530) );
  XNOR2_X1 U404 ( .A(n395), .B(KEYINPUT0), .ZN(n533) );
  AND2_X1 U405 ( .A1(G953), .A2(G902), .ZN(n479) );
  XNOR2_X1 U406 ( .A(n445), .B(n413), .ZN(n728) );
  XNOR2_X1 U407 ( .A(n446), .B(G134), .ZN(n413) );
  XNOR2_X1 U408 ( .A(G116), .B(G107), .ZN(n426) );
  NOR2_X1 U409 ( .A1(n555), .A2(n572), .ZN(n365) );
  NOR2_X1 U410 ( .A1(n543), .A2(n738), .ZN(n544) );
  XNOR2_X1 U411 ( .A(n728), .B(n447), .ZN(n524) );
  INV_X1 U412 ( .A(G146), .ZN(n447) );
  XNOR2_X1 U413 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n455) );
  OR2_X1 U414 ( .A1(n618), .A2(n617), .ZN(n619) );
  INV_X1 U415 ( .A(n375), .ZN(n723) );
  XNOR2_X1 U416 ( .A(n506), .B(n462), .ZN(n729) );
  XNOR2_X1 U417 ( .A(n456), .B(n417), .ZN(n458) );
  INV_X1 U418 ( .A(KEYINPUT23), .ZN(n417) );
  NAND2_X1 U419 ( .A1(G234), .A2(n731), .ZN(n463) );
  XOR2_X1 U420 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n464) );
  XNOR2_X1 U421 ( .A(n460), .B(n459), .ZN(n506) );
  INV_X1 U422 ( .A(KEYINPUT10), .ZN(n459) );
  OR2_X1 U423 ( .A1(n617), .A2(n471), .ZN(n397) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n371) );
  INV_X1 U425 ( .A(KEYINPUT83), .ZN(n358) );
  AND2_X1 U426 ( .A1(n601), .A2(n360), .ZN(n590) );
  AND2_X1 U427 ( .A1(n602), .A2(n653), .ZN(n360) );
  NAND2_X1 U428 ( .A1(n599), .A2(n384), .ZN(n383) );
  NOR2_X1 U429 ( .A1(n692), .A2(n533), .ZN(n536) );
  OR2_X1 U430 ( .A1(n548), .A2(n549), .ZN(n593) );
  XNOR2_X1 U431 ( .A(n403), .B(KEYINPUT107), .ZN(n402) );
  XNOR2_X1 U432 ( .A(n547), .B(n387), .ZN(n549) );
  INV_X1 U433 ( .A(KEYINPUT97), .ZN(n387) );
  XNOR2_X1 U434 ( .A(n396), .B(KEYINPUT19), .ZN(n571) );
  XNOR2_X1 U435 ( .A(n378), .B(KEYINPUT109), .ZN(n584) );
  XNOR2_X1 U436 ( .A(n363), .B(n362), .ZN(n570) );
  NOR2_X1 U437 ( .A1(n533), .A2(n512), .ZN(n513) );
  XNOR2_X1 U438 ( .A(n466), .B(n467), .ZN(n485) );
  XOR2_X1 U439 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n467) );
  XOR2_X1 U440 ( .A(KEYINPUT73), .B(KEYINPUT93), .Z(n516) );
  XNOR2_X1 U441 ( .A(G137), .B(G119), .ZN(n517) );
  XOR2_X1 U442 ( .A(KEYINPUT5), .B(G116), .Z(n518) );
  INV_X1 U443 ( .A(G125), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U445 ( .A(G110), .B(G101), .ZN(n448) );
  XOR2_X1 U446 ( .A(G107), .B(G104), .Z(n449) );
  XOR2_X1 U447 ( .A(G137), .B(G140), .Z(n461) );
  INV_X1 U448 ( .A(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U449 ( .A(KEYINPUT86), .B(KEYINPUT74), .ZN(n435) );
  NAND2_X1 U450 ( .A1(G237), .A2(G234), .ZN(n477) );
  OR2_X1 U451 ( .A1(n617), .A2(n420), .ZN(n419) );
  INV_X1 U452 ( .A(KEYINPUT2), .ZN(n420) );
  XNOR2_X1 U453 ( .A(n566), .B(KEYINPUT67), .ZN(n596) );
  INV_X1 U454 ( .A(KEYINPUT38), .ZN(n405) );
  XNOR2_X1 U455 ( .A(n510), .B(n509), .ZN(n547) );
  XNOR2_X1 U456 ( .A(n406), .B(n475), .ZN(n598) );
  XNOR2_X1 U457 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U458 ( .A(KEYINPUT28), .ZN(n362) );
  NAND2_X1 U459 ( .A1(n666), .A2(n665), .ZN(n671) );
  BUF_X1 U460 ( .A(n585), .Z(n567) );
  INV_X1 U461 ( .A(n562), .ZN(n665) );
  XOR2_X1 U462 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n493) );
  INV_X1 U463 ( .A(KEYINPUT95), .ZN(n392) );
  XNOR2_X1 U464 ( .A(n505), .B(n504), .ZN(n389) );
  XNOR2_X1 U465 ( .A(G140), .B(G113), .ZN(n501) );
  XOR2_X1 U466 ( .A(G131), .B(G143), .Z(n502) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n692) );
  INV_X1 U468 ( .A(KEYINPUT33), .ZN(n411) );
  NOR2_X1 U469 ( .A1(n723), .A2(n619), .ZN(n688) );
  NOR2_X1 U470 ( .A1(n671), .A2(n568), .ZN(n589) );
  XNOR2_X1 U471 ( .A(n398), .B(n352), .ZN(n714) );
  XNOR2_X1 U472 ( .A(n729), .B(n465), .ZN(n398) );
  XNOR2_X1 U473 ( .A(G128), .B(KEYINPUT24), .ZN(n457) );
  XNOR2_X1 U474 ( .A(n390), .B(n388), .ZN(n705) );
  XNOR2_X1 U475 ( .A(n507), .B(n391), .ZN(n390) );
  XNOR2_X1 U476 ( .A(n506), .B(n389), .ZN(n388) );
  XNOR2_X1 U477 ( .A(n503), .B(n392), .ZN(n391) );
  NAND2_X1 U478 ( .A1(n373), .A2(n620), .ZN(n372) );
  NOR2_X1 U479 ( .A1(G952), .A2(n731), .ZN(n717) );
  XNOR2_X1 U480 ( .A(n408), .B(n407), .ZN(n745) );
  INV_X1 U481 ( .A(KEYINPUT42), .ZN(n407) );
  XNOR2_X1 U482 ( .A(n591), .B(KEYINPUT40), .ZN(n743) );
  AND2_X1 U483 ( .A1(n380), .A2(n383), .ZN(n382) );
  XNOR2_X1 U484 ( .A(n542), .B(n541), .ZN(n738) );
  NOR2_X1 U485 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U486 ( .A(n368), .B(n367), .ZN(n742) );
  INV_X1 U487 ( .A(KEYINPUT32), .ZN(n367) );
  NOR2_X1 U488 ( .A1(n533), .A2(n677), .ZN(n552) );
  XNOR2_X1 U489 ( .A(n593), .B(n386), .ZN(n644) );
  INV_X1 U490 ( .A(KEYINPUT103), .ZN(n386) );
  AND2_X1 U491 ( .A1(n402), .A2(n401), .ZN(n605) );
  INV_X1 U492 ( .A(KEYINPUT77), .ZN(n376) );
  INV_X1 U493 ( .A(n594), .ZN(n393) );
  XNOR2_X1 U494 ( .A(n697), .B(n364), .ZN(G75) );
  XNOR2_X1 U495 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n364) );
  XNOR2_X1 U496 ( .A(n458), .B(n457), .ZN(n352) );
  XOR2_X1 U497 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n353) );
  XOR2_X1 U498 ( .A(KEYINPUT101), .B(n556), .Z(n354) );
  AND2_X1 U499 ( .A1(n607), .A2(KEYINPUT79), .ZN(n355) );
  AND2_X1 U500 ( .A1(n614), .A2(KEYINPUT36), .ZN(n356) );
  XNOR2_X1 U501 ( .A(G902), .B(KEYINPUT15), .ZN(n471) );
  NOR2_X1 U502 ( .A1(n421), .A2(n423), .ZN(n357) );
  NOR2_X1 U503 ( .A1(n743), .A2(n745), .ZN(n422) );
  XNOR2_X2 U504 ( .A(n361), .B(n609), .ZN(n618) );
  NAND2_X1 U505 ( .A1(n596), .A2(n567), .ZN(n363) );
  INV_X1 U506 ( .A(n400), .ZN(n690) );
  NAND2_X1 U507 ( .A1(n485), .A2(G221), .ZN(n486) );
  NAND2_X1 U508 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X2 U509 ( .A(n410), .B(KEYINPUT45), .ZN(n375) );
  BUF_X2 U510 ( .A(n598), .Z(n614) );
  INV_X1 U511 ( .A(n426), .ZN(n490) );
  XOR2_X1 U512 ( .A(n452), .B(n451), .Z(n453) );
  XNOR2_X1 U513 ( .A(n524), .B(n453), .ZN(n698) );
  NOR2_X1 U514 ( .A1(n365), .A2(n632), .ZN(n556) );
  XNOR2_X1 U515 ( .A(n366), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U516 ( .A(n430), .B(n431), .ZN(n434) );
  NAND2_X1 U517 ( .A1(n530), .A2(n529), .ZN(n368) );
  XNOR2_X1 U518 ( .A(n369), .B(KEYINPUT126), .ZN(G66) );
  NOR2_X2 U519 ( .A1(n716), .A2(n717), .ZN(n369) );
  NOR2_X1 U520 ( .A1(n618), .A2(n397), .ZN(n374) );
  XNOR2_X2 U521 ( .A(n377), .B(n376), .ZN(n643) );
  NAND2_X1 U522 ( .A1(n584), .A2(n571), .ZN(n377) );
  NAND2_X1 U523 ( .A1(n570), .A2(n569), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n379), .A2(n356), .ZN(n381) );
  INV_X1 U525 ( .A(n610), .ZN(n379) );
  NAND2_X1 U526 ( .A1(n610), .A2(n384), .ZN(n380) );
  NAND2_X1 U527 ( .A1(n382), .A2(n381), .ZN(n385) );
  INV_X1 U528 ( .A(KEYINPUT36), .ZN(n384) );
  NAND2_X1 U529 ( .A1(n385), .A2(n611), .ZN(n600) );
  INV_X1 U530 ( .A(n644), .ZN(n646) );
  AND2_X1 U531 ( .A1(n394), .A2(n393), .ZN(n545) );
  XNOR2_X1 U532 ( .A(n513), .B(KEYINPUT22), .ZN(n394) );
  NAND2_X1 U533 ( .A1(n571), .A2(n484), .ZN(n395) );
  NAND2_X1 U534 ( .A1(n598), .A2(n654), .ZN(n396) );
  INV_X1 U535 ( .A(n603), .ZN(n401) );
  NAND2_X1 U536 ( .A1(n601), .A2(n404), .ZN(n403) );
  AND2_X1 U537 ( .A1(n602), .A2(n614), .ZN(n404) );
  NAND2_X1 U538 ( .A1(n653), .A2(n654), .ZN(n582) );
  NAND2_X1 U539 ( .A1(n472), .A2(n471), .ZN(n406) );
  NAND2_X1 U540 ( .A1(n679), .A2(n584), .ZN(n408) );
  NAND2_X1 U541 ( .A1(n354), .A2(n409), .ZN(n410) );
  XNOR2_X1 U542 ( .A(n544), .B(KEYINPUT44), .ZN(n409) );
  NAND2_X1 U543 ( .A1(n550), .A2(n594), .ZN(n412) );
  XNOR2_X1 U544 ( .A(n534), .B(KEYINPUT72), .ZN(n550) );
  XNOR2_X1 U545 ( .A(n619), .B(n730), .ZN(n732) );
  XNOR2_X1 U546 ( .A(n422), .B(n592), .ZN(n421) );
  NAND2_X1 U547 ( .A1(n425), .A2(n424), .ZN(n423) );
  NOR2_X1 U548 ( .A1(n739), .A2(n355), .ZN(n424) );
  INV_X1 U549 ( .A(n606), .ZN(n425) );
  INV_X1 U550 ( .A(KEYINPUT46), .ZN(n592) );
  XNOR2_X1 U551 ( .A(n445), .B(n438), .ZN(n439) );
  INV_X1 U552 ( .A(n461), .ZN(n462) );
  XNOR2_X1 U553 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n522), .B(n433), .ZN(n523) );
  XNOR2_X1 U555 ( .A(n524), .B(n523), .ZN(n625) );
  XNOR2_X1 U556 ( .A(n705), .B(n704), .ZN(n706) );
  INV_X1 U557 ( .A(KEYINPUT35), .ZN(n541) );
  XNOR2_X1 U558 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n443) );
  NAND2_X1 U559 ( .A1(KEYINPUT16), .A2(n426), .ZN(n429) );
  INV_X1 U560 ( .A(KEYINPUT16), .ZN(n427) );
  NAND2_X1 U561 ( .A1(n427), .A2(n490), .ZN(n428) );
  NAND2_X1 U562 ( .A1(n429), .A2(n428), .ZN(n431) );
  XNOR2_X1 U563 ( .A(n505), .B(n456), .ZN(n430) );
  XOR2_X1 U564 ( .A(G101), .B(KEYINPUT3), .Z(n432) );
  XOR2_X1 U565 ( .A(G113), .B(n432), .Z(n433) );
  INV_X1 U566 ( .A(n433), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n434), .B(n521), .ZN(n718) );
  XNOR2_X1 U568 ( .A(n353), .B(n435), .ZN(n437) );
  INV_X1 U569 ( .A(n460), .ZN(n436) );
  XNOR2_X1 U570 ( .A(n437), .B(n436), .ZN(n440) );
  NAND2_X1 U571 ( .A1(G224), .A2(n731), .ZN(n438) );
  XNOR2_X1 U572 ( .A(n718), .B(n441), .ZN(n472) );
  XNOR2_X1 U573 ( .A(n472), .B(KEYINPUT122), .ZN(n442) );
  XNOR2_X1 U574 ( .A(n443), .B(n442), .ZN(n622) );
  XOR2_X1 U575 ( .A(n471), .B(KEYINPUT82), .Z(n444) );
  NAND2_X1 U576 ( .A1(n444), .A2(KEYINPUT2), .ZN(n620) );
  INV_X1 U577 ( .A(G131), .ZN(n446) );
  XOR2_X1 U578 ( .A(n461), .B(n450), .Z(n452) );
  NAND2_X1 U579 ( .A1(G227), .A2(n731), .ZN(n451) );
  INV_X1 U580 ( .A(n670), .ZN(n611) );
  XNOR2_X1 U581 ( .A(n464), .B(n463), .ZN(n496) );
  NAND2_X1 U582 ( .A1(G221), .A2(n496), .ZN(n465) );
  XOR2_X1 U583 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n469) );
  NAND2_X1 U584 ( .A1(G234), .A2(n471), .ZN(n466) );
  NAND2_X1 U585 ( .A1(n485), .A2(G217), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U587 ( .A1(G210), .A2(n476), .ZN(n474) );
  INV_X1 U588 ( .A(KEYINPUT78), .ZN(n473) );
  NAND2_X1 U589 ( .A1(G214), .A2(n476), .ZN(n654) );
  XNOR2_X1 U590 ( .A(n477), .B(KEYINPUT14), .ZN(n480) );
  NAND2_X1 U591 ( .A1(n480), .A2(G952), .ZN(n478) );
  XOR2_X1 U592 ( .A(KEYINPUT87), .B(n478), .Z(n685) );
  NOR2_X1 U593 ( .A1(G953), .A2(n685), .ZN(n561) );
  NAND2_X1 U594 ( .A1(n480), .A2(n479), .ZN(n557) );
  NOR2_X1 U595 ( .A1(G898), .A2(n557), .ZN(n481) );
  XNOR2_X1 U596 ( .A(n481), .B(KEYINPUT88), .ZN(n482) );
  NOR2_X1 U597 ( .A1(n561), .A2(n482), .ZN(n483) );
  XNOR2_X1 U598 ( .A(KEYINPUT89), .B(n483), .ZN(n484) );
  XNOR2_X1 U599 ( .A(n486), .B(KEYINPUT92), .ZN(n487) );
  XNOR2_X1 U600 ( .A(KEYINPUT100), .B(G478), .ZN(n500) );
  XOR2_X1 U601 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n489) );
  XNOR2_X1 U602 ( .A(G122), .B(G134), .ZN(n488) );
  XNOR2_X1 U603 ( .A(n489), .B(n488), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U606 ( .A(n495), .B(n494), .Z(n498) );
  NAND2_X1 U607 ( .A1(G217), .A2(n496), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n498), .B(n497), .ZN(n709) );
  NOR2_X1 U609 ( .A1(G902), .A2(n709), .ZN(n499) );
  XOR2_X1 U610 ( .A(n500), .B(n499), .Z(n548) );
  INV_X1 U611 ( .A(n548), .ZN(n537) );
  XNOR2_X1 U612 ( .A(n502), .B(n501), .ZN(n507) );
  XOR2_X1 U613 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n504) );
  NAND2_X1 U614 ( .A1(n514), .A2(G214), .ZN(n503) );
  NOR2_X1 U615 ( .A1(n705), .A2(G902), .ZN(n510) );
  XOR2_X1 U616 ( .A(G475), .B(KEYINPUT13), .Z(n508) );
  XNOR2_X1 U617 ( .A(KEYINPUT96), .B(n508), .ZN(n509) );
  NAND2_X1 U618 ( .A1(n537), .A2(n547), .ZN(n657) );
  INV_X1 U619 ( .A(n657), .ZN(n511) );
  NAND2_X1 U620 ( .A1(n665), .A2(n511), .ZN(n512) );
  NAND2_X1 U621 ( .A1(n514), .A2(G210), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U624 ( .A(n520), .B(n519), .Z(n522) );
  NOR2_X1 U625 ( .A1(n625), .A2(G902), .ZN(n526) );
  INV_X1 U626 ( .A(G472), .ZN(n525) );
  INV_X1 U627 ( .A(n567), .ZN(n553) );
  NAND2_X1 U628 ( .A1(n530), .A2(n553), .ZN(n527) );
  NOR2_X1 U629 ( .A1(n611), .A2(n527), .ZN(n639) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n585), .Z(n594) );
  XOR2_X1 U631 ( .A(KEYINPUT76), .B(n594), .Z(n528) );
  AND2_X1 U632 ( .A1(n528), .A2(n611), .ZN(n529) );
  NOR2_X1 U633 ( .A1(n639), .A2(n742), .ZN(n532) );
  INV_X1 U634 ( .A(KEYINPUT84), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n543) );
  NOR2_X1 U636 ( .A1(n670), .A2(n671), .ZN(n534) );
  XNOR2_X1 U637 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n535) );
  XNOR2_X1 U638 ( .A(n536), .B(n535), .ZN(n540) );
  NOR2_X1 U639 ( .A1(n537), .A2(n547), .ZN(n538) );
  XOR2_X1 U640 ( .A(KEYINPUT102), .B(n538), .Z(n603) );
  XOR2_X1 U641 ( .A(n603), .B(KEYINPUT75), .Z(n539) );
  NAND2_X1 U642 ( .A1(n666), .A2(n545), .ZN(n546) );
  NOR2_X1 U643 ( .A1(n611), .A2(n546), .ZN(n632) );
  NAND2_X1 U644 ( .A1(n549), .A2(n548), .ZN(n640) );
  NAND2_X1 U645 ( .A1(n593), .A2(n640), .ZN(n576) );
  INV_X1 U646 ( .A(n576), .ZN(n660) );
  XNOR2_X1 U647 ( .A(KEYINPUT80), .B(n660), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n550), .A2(n567), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n551), .B(KEYINPUT94), .ZN(n677) );
  XOR2_X1 U650 ( .A(KEYINPUT31), .B(n552), .Z(n649) );
  NAND2_X1 U651 ( .A1(n589), .A2(n553), .ZN(n554) );
  NOR2_X1 U652 ( .A1(n533), .A2(n554), .ZN(n635) );
  NOR2_X1 U653 ( .A1(n649), .A2(n635), .ZN(n555) );
  XNOR2_X1 U654 ( .A(KEYINPUT104), .B(n557), .ZN(n558) );
  NOR2_X1 U655 ( .A1(G900), .A2(n558), .ZN(n559) );
  XOR2_X1 U656 ( .A(KEYINPUT105), .B(n559), .Z(n560) );
  NOR2_X1 U657 ( .A1(n561), .A2(n560), .ZN(n588) );
  NOR2_X1 U658 ( .A1(n588), .A2(n562), .ZN(n563) );
  XNOR2_X1 U659 ( .A(n563), .B(KEYINPUT68), .ZN(n565) );
  INV_X1 U660 ( .A(n666), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U662 ( .A(n568), .ZN(n569) );
  NOR2_X1 U663 ( .A1(KEYINPUT47), .A2(n572), .ZN(n573) );
  XNOR2_X1 U664 ( .A(KEYINPUT71), .B(n573), .ZN(n574) );
  XNOR2_X1 U665 ( .A(KEYINPUT70), .B(n575), .ZN(n581) );
  INV_X1 U666 ( .A(KEYINPUT47), .ZN(n579) );
  NOR2_X1 U667 ( .A1(KEYINPUT79), .A2(n576), .ZN(n577) );
  NOR2_X1 U668 ( .A1(n643), .A2(n577), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U670 ( .A1(n581), .A2(n580), .ZN(n608) );
  XNOR2_X1 U671 ( .A(n582), .B(KEYINPUT110), .ZN(n659) );
  XNOR2_X1 U672 ( .A(n583), .B(KEYINPUT41), .ZN(n691) );
  NAND2_X1 U673 ( .A1(n585), .A2(n654), .ZN(n586) );
  XNOR2_X1 U674 ( .A(KEYINPUT30), .B(n586), .ZN(n587) );
  NOR2_X1 U675 ( .A1(n588), .A2(n587), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n589), .B(KEYINPUT106), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n590), .B(KEYINPUT39), .ZN(n615) );
  NOR2_X1 U678 ( .A1(n615), .A2(n593), .ZN(n591) );
  NAND2_X1 U679 ( .A1(n594), .A2(n654), .ZN(n595) );
  NOR2_X1 U680 ( .A1(n644), .A2(n595), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n610) );
  INV_X1 U682 ( .A(n614), .ZN(n599) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT111), .ZN(n739) );
  INV_X1 U684 ( .A(KEYINPUT108), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n605), .B(n604), .ZN(n744) );
  XNOR2_X1 U686 ( .A(n744), .B(KEYINPUT81), .ZN(n606) );
  NAND2_X1 U687 ( .A1(KEYINPUT47), .A2(n660), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n652) );
  OR2_X1 U691 ( .A1(n615), .A2(n640), .ZN(n651) );
  NAND2_X1 U692 ( .A1(n710), .A2(G210), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X2 U694 ( .A1(n623), .A2(n717), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U696 ( .A1(n710), .A2(G472), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT62), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(KEYINPUT85), .B(KEYINPUT112), .ZN(n629) );
  XNOR2_X1 U700 ( .A(n629), .B(KEYINPUT63), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(G57) );
  XOR2_X1 U702 ( .A(G101), .B(n632), .Z(G3) );
  XOR2_X1 U703 ( .A(G104), .B(KEYINPUT113), .Z(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n646), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  INV_X1 U707 ( .A(n640), .ZN(n648) );
  NAND2_X1 U708 ( .A1(n635), .A2(n648), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U710 ( .A(G107), .B(n638), .ZN(G9) );
  XOR2_X1 U711 ( .A(G110), .B(n639), .Z(G12) );
  NOR2_X1 U712 ( .A1(n640), .A2(n643), .ZN(n642) );
  XNOR2_X1 U713 ( .A(G128), .B(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(G30) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U716 ( .A(G146), .B(n645), .Z(G48) );
  NAND2_X1 U717 ( .A1(n649), .A2(n646), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(G113), .ZN(G15) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(G116), .ZN(G18) );
  XNOR2_X1 U721 ( .A(G134), .B(n651), .ZN(G36) );
  XOR2_X1 U722 ( .A(G140), .B(n652), .Z(G42) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U724 ( .A(KEYINPUT117), .B(n655), .Z(n656) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT118), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U729 ( .A1(n663), .A2(n692), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(KEYINPUT119), .ZN(n682) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT49), .B(n667), .Z(n668) );
  NOR2_X1 U733 ( .A1(n567), .A2(n668), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT115), .B(n669), .Z(n675) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n672), .B(KEYINPUT116), .ZN(n673) );
  XNOR2_X1 U737 ( .A(KEYINPUT50), .B(n673), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n678), .Z(n680) );
  NAND2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n684) );
  XOR2_X1 U743 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n683) );
  XNOR2_X1 U744 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U746 ( .A1(G953), .A2(n687), .ZN(n696) );
  NOR2_X1 U747 ( .A1(KEYINPUT2), .A2(n688), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U751 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT123), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U755 ( .A1(n710), .A2(G469), .ZN(n701) );
  XOR2_X1 U756 ( .A(n702), .B(n701), .Z(n703) );
  NOR2_X1 U757 ( .A1(n717), .A2(n703), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n710), .A2(G475), .ZN(n707) );
  XOR2_X1 U759 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n704) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  XOR2_X1 U761 ( .A(n709), .B(KEYINPUT125), .Z(n712) );
  NAND2_X1 U762 ( .A1(n710), .A2(G478), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n717), .A2(n713), .ZN(G63) );
  NAND2_X1 U765 ( .A1(G217), .A2(n710), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  OR2_X1 U767 ( .A1(G898), .A2(n731), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n727) );
  NAND2_X1 U769 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U771 ( .A1(n721), .A2(G898), .ZN(n722) );
  XNOR2_X1 U772 ( .A(n722), .B(KEYINPUT127), .ZN(n725) );
  NOR2_X1 U773 ( .A1(n723), .A2(G953), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U776 ( .A(n729), .B(n728), .ZN(n733) );
  INV_X1 U777 ( .A(n733), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n732), .A2(n731), .ZN(n737) );
  XOR2_X1 U779 ( .A(G227), .B(n733), .Z(n734) );
  NAND2_X1 U780 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U783 ( .A(n738), .B(G122), .Z(G24) );
  XNOR2_X1 U784 ( .A(n739), .B(KEYINPUT37), .ZN(n740) );
  XNOR2_X1 U785 ( .A(n740), .B(KEYINPUT114), .ZN(n741) );
  XNOR2_X1 U786 ( .A(G125), .B(n741), .ZN(G27) );
  XOR2_X1 U787 ( .A(n742), .B(G119), .Z(G21) );
  XOR2_X1 U788 ( .A(n743), .B(G131), .Z(G33) );
  XNOR2_X1 U789 ( .A(n744), .B(G143), .ZN(G45) );
  XOR2_X1 U790 ( .A(n745), .B(G137), .Z(G39) );
endmodule

