

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746;

  NAND2_X1 U369 ( .A1(n387), .A2(n391), .ZN(n576) );
  INV_X1 U370 ( .A(n509), .ZN(n484) );
  NAND2_X1 U371 ( .A1(n588), .A2(n581), .ZN(n573) );
  NOR2_X1 U372 ( .A1(n564), .A2(n670), .ZN(n499) );
  NAND2_X1 U373 ( .A1(n384), .A2(n381), .ZN(n534) );
  XNOR2_X1 U374 ( .A(n505), .B(n504), .ZN(n712) );
  XNOR2_X1 U375 ( .A(n725), .B(KEYINPUT72), .ZN(n503) );
  XNOR2_X1 U376 ( .A(n394), .B(G101), .ZN(n393) );
  BUF_X1 U377 ( .A(G113), .Z(n348) );
  AND2_X2 U378 ( .A1(n666), .A2(n665), .ZN(n588) );
  XNOR2_X2 U379 ( .A(n478), .B(G122), .ZN(n423) );
  INV_X1 U380 ( .A(n348), .ZN(n445) );
  INV_X1 U381 ( .A(G953), .ZN(n736) );
  NAND2_X2 U382 ( .A1(n570), .A2(n569), .ZN(n577) );
  NAND2_X2 U383 ( .A1(n403), .A2(n401), .ZN(n596) );
  AND2_X2 U384 ( .A1(n404), .A2(n595), .ZN(n403) );
  XNOR2_X2 U385 ( .A(n734), .B(G146), .ZN(n505) );
  XNOR2_X2 U386 ( .A(n576), .B(KEYINPUT35), .ZN(n627) );
  XNOR2_X1 U387 ( .A(n418), .B(n416), .ZN(n744) );
  XNOR2_X1 U388 ( .A(n509), .B(KEYINPUT6), .ZN(n581) );
  XNOR2_X1 U389 ( .A(n619), .B(n618), .ZN(n620) );
  OR2_X1 U390 ( .A1(n717), .A2(G902), .ZN(n495) );
  XNOR2_X1 U391 ( .A(G137), .B(G134), .ZN(n470) );
  XNOR2_X2 U392 ( .A(n423), .B(n424), .ZN(n726) );
  XNOR2_X2 U393 ( .A(n409), .B(n408), .ZN(n725) );
  XNOR2_X2 U394 ( .A(G110), .B(G107), .ZN(n409) );
  XNOR2_X1 U395 ( .A(KEYINPUT68), .B(G131), .ZN(n471) );
  XNOR2_X1 U396 ( .A(n443), .B(n444), .ZN(n732) );
  XOR2_X1 U397 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n444) );
  XNOR2_X1 U398 ( .A(n522), .B(KEYINPUT39), .ZN(n541) );
  XNOR2_X1 U399 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n561) );
  XNOR2_X1 U400 ( .A(n493), .B(KEYINPUT25), .ZN(n494) );
  NAND2_X1 U401 ( .A1(n506), .A2(G902), .ZN(n385) );
  AND2_X1 U402 ( .A1(n539), .A2(n352), .ZN(n368) );
  NAND2_X1 U403 ( .A1(n579), .A2(n578), .ZN(n402) );
  OR2_X1 U404 ( .A1(n627), .A2(KEYINPUT44), .ZN(n579) );
  INV_X1 U405 ( .A(G128), .ZN(n425) );
  XNOR2_X1 U406 ( .A(G143), .B(G104), .ZN(n438) );
  XNOR2_X1 U407 ( .A(n534), .B(KEYINPUT1), .ZN(n565) );
  XNOR2_X1 U408 ( .A(n375), .B(n356), .ZN(n697) );
  NOR2_X1 U409 ( .A1(n682), .A2(n377), .ZN(n376) );
  INV_X1 U410 ( .A(n523), .ZN(n530) );
  BUF_X1 U411 ( .A(n565), .Z(n369) );
  AND2_X1 U412 ( .A1(n581), .A2(n354), .ZN(n398) );
  NOR2_X1 U413 ( .A1(n413), .A2(n415), .ZN(n507) );
  XNOR2_X1 U414 ( .A(n485), .B(KEYINPUT30), .ZN(n415) );
  XNOR2_X1 U415 ( .A(n450), .B(n628), .ZN(n524) );
  NOR2_X1 U416 ( .A1(n364), .A2(n719), .ZN(n363) );
  NOR2_X1 U417 ( .A1(n367), .A2(G472), .ZN(n364) );
  NAND2_X1 U418 ( .A1(n362), .A2(n625), .ZN(n361) );
  INV_X1 U419 ( .A(G217), .ZN(n422) );
  XNOR2_X1 U420 ( .A(n373), .B(n489), .ZN(n717) );
  XNOR2_X1 U421 ( .A(n732), .B(n491), .ZN(n373) );
  XOR2_X1 U422 ( .A(G119), .B(G137), .Z(n487) );
  INV_X1 U423 ( .A(KEYINPUT124), .ZN(n420) );
  XNOR2_X1 U424 ( .A(n480), .B(KEYINPUT15), .ZN(n601) );
  XNOR2_X1 U425 ( .A(n428), .B(G146), .ZN(n442) );
  INV_X1 U426 ( .A(G125), .ZN(n428) );
  XNOR2_X1 U427 ( .A(G107), .B(G134), .ZN(n451) );
  XNOR2_X1 U428 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U429 ( .A(n379), .B(n378), .ZN(n431) );
  XNOR2_X1 U430 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n380), .B(KEYINPUT88), .ZN(n379) );
  XNOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n380) );
  INV_X1 U433 ( .A(n679), .ZN(n377) );
  INV_X1 U434 ( .A(n565), .ZN(n665) );
  XNOR2_X1 U435 ( .A(n505), .B(n479), .ZN(n624) );
  AND2_X1 U436 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U437 ( .A1(n383), .A2(n480), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n540), .B(KEYINPUT48), .ZN(n549) );
  INV_X1 U439 ( .A(G104), .ZN(n408) );
  XNOR2_X1 U440 ( .A(n372), .B(n350), .ZN(n488) );
  XNOR2_X1 U441 ( .A(n486), .B(KEYINPUT23), .ZN(n372) );
  XNOR2_X1 U442 ( .A(G128), .B(G110), .ZN(n486) );
  XNOR2_X1 U443 ( .A(n399), .B(n732), .ZN(n630) );
  XNOR2_X1 U444 ( .A(n447), .B(n400), .ZN(n399) );
  XNOR2_X1 U445 ( .A(n446), .B(G122), .ZN(n400) );
  XOR2_X1 U446 ( .A(G140), .B(G101), .Z(n501) );
  NAND2_X1 U447 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U448 ( .A(n610), .ZN(n611) );
  NOR2_X1 U449 ( .A1(n697), .A2(n526), .ZN(n528) );
  XNOR2_X1 U450 ( .A(n417), .B(KEYINPUT40), .ZN(n416) );
  NAND2_X1 U451 ( .A1(n541), .A2(n530), .ZN(n418) );
  INV_X1 U452 ( .A(KEYINPUT105), .ZN(n417) );
  NOR2_X1 U453 ( .A1(n545), .A2(n349), .ZN(n533) );
  XNOR2_X1 U454 ( .A(n410), .B(n568), .ZN(n743) );
  AND2_X1 U455 ( .A1(n567), .A2(n412), .ZN(n411) );
  XNOR2_X1 U456 ( .A(n523), .B(KEYINPUT103), .ZN(n652) );
  XNOR2_X1 U457 ( .A(n366), .B(n359), .ZN(G57) );
  NAND2_X1 U458 ( .A1(n351), .A2(n361), .ZN(n366) );
  XNOR2_X1 U459 ( .A(n421), .B(n419), .ZN(n718) );
  XNOR2_X1 U460 ( .A(n717), .B(n420), .ZN(n419) );
  NOR2_X1 U461 ( .A1(n362), .A2(n422), .ZN(n421) );
  NAND2_X1 U462 ( .A1(n652), .A2(n398), .ZN(n349) );
  XOR2_X1 U463 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n350) );
  AND2_X1 U464 ( .A1(n365), .A2(n363), .ZN(n351) );
  XOR2_X1 U465 ( .A(KEYINPUT82), .B(n521), .Z(n352) );
  XOR2_X1 U466 ( .A(n529), .B(KEYINPUT46), .Z(n353) );
  AND2_X1 U467 ( .A1(n532), .A2(n679), .ZN(n354) );
  OR2_X1 U468 ( .A1(n586), .A2(KEYINPUT34), .ZN(n355) );
  XOR2_X1 U469 ( .A(KEYINPUT41), .B(KEYINPUT106), .Z(n356) );
  AND2_X1 U470 ( .A1(n367), .A2(G472), .ZN(n357) );
  OR2_X1 U471 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n358) );
  INV_X1 U472 ( .A(n625), .ZN(n367) );
  XOR2_X1 U473 ( .A(KEYINPUT62), .B(n624), .Z(n625) );
  XOR2_X1 U474 ( .A(KEYINPUT63), .B(KEYINPUT109), .Z(n359) );
  NAND2_X1 U475 ( .A1(n360), .A2(n411), .ZN(n410) );
  AND2_X2 U476 ( .A1(n360), .A2(n369), .ZN(n583) );
  XNOR2_X2 U477 ( .A(n562), .B(n561), .ZN(n360) );
  INV_X1 U478 ( .A(n716), .ZN(n362) );
  NAND2_X1 U479 ( .A1(n716), .A2(n357), .ZN(n365) );
  NAND2_X1 U480 ( .A1(n368), .A2(n353), .ZN(n540) );
  OR2_X1 U481 ( .A1(n535), .A2(n369), .ZN(n661) );
  XNOR2_X2 U482 ( .A(n482), .B(n481), .ZN(n509) );
  NAND2_X2 U483 ( .A1(n370), .A2(n704), .ZN(n629) );
  NAND2_X1 U484 ( .A1(n604), .A2(n605), .ZN(n370) );
  XNOR2_X1 U485 ( .A(n371), .B(n726), .ZN(n617) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n371) );
  XNOR2_X1 U487 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U488 ( .A(n629), .ZN(n716) );
  NAND2_X1 U489 ( .A1(n374), .A2(n563), .ZN(n570) );
  XNOR2_X1 U490 ( .A(n583), .B(KEYINPUT102), .ZN(n374) );
  NOR2_X2 U491 ( .A1(n549), .A2(n548), .ZN(n735) );
  NOR2_X2 U492 ( .A1(n545), .A2(n508), .ZN(n650) );
  NAND2_X1 U493 ( .A1(n376), .A2(n680), .ZN(n375) );
  NAND2_X1 U494 ( .A1(n680), .A2(n679), .ZN(n685) );
  OR2_X1 U495 ( .A1(n712), .A2(n382), .ZN(n381) );
  INV_X1 U496 ( .A(n506), .ZN(n383) );
  NAND2_X1 U497 ( .A1(n712), .A2(n506), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U499 ( .A1(n698), .A2(n574), .ZN(n388) );
  NAND2_X1 U500 ( .A1(n390), .A2(n355), .ZN(n389) );
  INV_X1 U501 ( .A(n698), .ZN(n390) );
  AND2_X1 U502 ( .A1(n392), .A2(n575), .ZN(n391) );
  NAND2_X1 U503 ( .A1(n586), .A2(KEYINPUT34), .ZN(n392) );
  XNOR2_X2 U504 ( .A(n573), .B(n572), .ZN(n698) );
  XNOR2_X2 U505 ( .A(n395), .B(n393), .ZN(n478) );
  XNOR2_X2 U506 ( .A(G119), .B(KEYINPUT71), .ZN(n394) );
  XNOR2_X2 U507 ( .A(n396), .B(n397), .ZN(n395) );
  XNOR2_X2 U508 ( .A(G116), .B(G113), .ZN(n396) );
  XNOR2_X2 U509 ( .A(KEYINPUT3), .B(KEYINPUT70), .ZN(n397) );
  INV_X1 U510 ( .A(n570), .ZN(n645) );
  NAND2_X1 U511 ( .A1(n402), .A2(n580), .ZN(n401) );
  NAND2_X1 U512 ( .A1(n405), .A2(n358), .ZN(n404) );
  NAND2_X1 U513 ( .A1(n571), .A2(n406), .ZN(n405) );
  NOR2_X1 U514 ( .A1(n627), .A2(n407), .ZN(n406) );
  INV_X1 U515 ( .A(KEYINPUT44), .ZN(n407) );
  INV_X1 U516 ( .A(n581), .ZN(n412) );
  NAND2_X1 U517 ( .A1(n666), .A2(n414), .ZN(n413) );
  NOR2_X1 U518 ( .A1(n534), .A2(n510), .ZN(n414) );
  NOR2_X2 U519 ( .A1(n614), .A2(n719), .ZN(n616) );
  XNOR2_X2 U520 ( .A(n473), .B(n472), .ZN(n734) );
  XNOR2_X2 U521 ( .A(n458), .B(n427), .ZN(n473) );
  XNOR2_X2 U522 ( .A(n426), .B(n425), .ZN(n458) );
  INV_X1 U523 ( .A(n531), .ZN(n532) );
  AND2_X1 U524 ( .A1(n661), .A2(n538), .ZN(n539) );
  XNOR2_X1 U525 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U526 ( .A(n471), .B(n445), .ZN(n446) );
  INV_X1 U527 ( .A(KEYINPUT0), .ZN(n556) );
  INV_X1 U528 ( .A(KEYINPUT123), .ZN(n615) );
  XNOR2_X1 U529 ( .A(n616), .B(n615), .ZN(G63) );
  INV_X1 U530 ( .A(G902), .ZN(n480) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n424) );
  XNOR2_X2 U532 ( .A(KEYINPUT80), .B(G143), .ZN(n426) );
  XNOR2_X1 U533 ( .A(n473), .B(n503), .ZN(n433) );
  NAND2_X1 U534 ( .A1(G224), .A2(n736), .ZN(n429) );
  XNOR2_X1 U535 ( .A(n442), .B(n429), .ZN(n430) );
  NOR2_X1 U536 ( .A1(n601), .A2(n617), .ZN(n435) );
  OR2_X1 U537 ( .A1(G902), .A2(G237), .ZN(n483) );
  NAND2_X1 U538 ( .A1(n483), .A2(G210), .ZN(n434) );
  XNOR2_X1 U539 ( .A(n435), .B(n434), .ZN(n514) );
  INV_X1 U540 ( .A(n514), .ZN(n545) );
  XOR2_X1 U541 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n437) );
  NOR2_X1 U542 ( .A1(G953), .A2(G237), .ZN(n474) );
  NAND2_X1 U543 ( .A1(n474), .A2(G214), .ZN(n436) );
  XNOR2_X1 U544 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U545 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n439) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n441), .B(n440), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n442), .B(G140), .ZN(n443) );
  NOR2_X1 U549 ( .A1(G902), .A2(n630), .ZN(n449) );
  XNOR2_X1 U550 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n448) );
  XNOR2_X1 U551 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U552 ( .A(G475), .ZN(n628) );
  XOR2_X1 U553 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n452) );
  XNOR2_X1 U554 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U555 ( .A(n453), .B(KEYINPUT7), .Z(n455) );
  XNOR2_X1 U556 ( .A(G116), .B(G122), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n461) );
  XOR2_X1 U558 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n457) );
  NAND2_X1 U559 ( .A1(G234), .A2(n736), .ZN(n456) );
  XNOR2_X1 U560 ( .A(n457), .B(n456), .ZN(n490) );
  NAND2_X1 U561 ( .A1(G217), .A2(n490), .ZN(n459) );
  XNOR2_X1 U562 ( .A(n458), .B(n459), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n461), .B(n460), .ZN(n610) );
  NAND2_X1 U564 ( .A1(n610), .A2(n480), .ZN(n463) );
  XOR2_X1 U565 ( .A(G478), .B(KEYINPUT99), .Z(n462) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n525) );
  AND2_X1 U567 ( .A1(n524), .A2(n525), .ZN(n575) );
  NAND2_X1 U568 ( .A1(G237), .A2(G234), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n464), .B(KEYINPUT14), .ZN(n466) );
  NAND2_X1 U570 ( .A1(G902), .A2(n466), .ZN(n550) );
  NOR2_X1 U571 ( .A1(G900), .A2(n550), .ZN(n465) );
  NAND2_X1 U572 ( .A1(n465), .A2(G953), .ZN(n468) );
  NAND2_X1 U573 ( .A1(G952), .A2(n466), .ZN(n467) );
  XNOR2_X1 U574 ( .A(KEYINPUT89), .B(n467), .ZN(n695) );
  NAND2_X1 U575 ( .A1(n695), .A2(n736), .ZN(n553) );
  NAND2_X1 U576 ( .A1(n468), .A2(n553), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n469), .B(KEYINPUT81), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U579 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n476) );
  NAND2_X1 U580 ( .A1(G210), .A2(n474), .ZN(n475) );
  XNOR2_X1 U581 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U583 ( .A1(n624), .A2(n480), .ZN(n482) );
  XOR2_X1 U584 ( .A(KEYINPUT74), .B(G472), .Z(n481) );
  NAND2_X1 U585 ( .A1(G214), .A2(n483), .ZN(n679) );
  NAND2_X1 U586 ( .A1(n484), .A2(n679), .ZN(n485) );
  XNOR2_X1 U587 ( .A(n488), .B(n487), .ZN(n489) );
  AND2_X1 U588 ( .A1(G221), .A2(n490), .ZN(n491) );
  INV_X1 U589 ( .A(n601), .ZN(n599) );
  NAND2_X1 U590 ( .A1(n599), .A2(G234), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n492), .B(KEYINPUT20), .ZN(n496) );
  NAND2_X1 U592 ( .A1(G217), .A2(n496), .ZN(n493) );
  XNOR2_X2 U593 ( .A(n495), .B(n494), .ZN(n564) );
  XOR2_X1 U594 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n498) );
  NAND2_X1 U595 ( .A1(G221), .A2(n496), .ZN(n497) );
  XNOR2_X1 U596 ( .A(n498), .B(n497), .ZN(n670) );
  XNOR2_X2 U597 ( .A(n499), .B(KEYINPUT66), .ZN(n666) );
  NAND2_X1 U598 ( .A1(G227), .A2(n736), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U601 ( .A(KEYINPUT69), .B(G469), .ZN(n506) );
  NAND2_X1 U602 ( .A1(n575), .A2(n507), .ZN(n508) );
  XNOR2_X1 U603 ( .A(n650), .B(KEYINPUT83), .ZN(n520) );
  NOR2_X1 U604 ( .A1(n670), .A2(n510), .ZN(n511) );
  NAND2_X1 U605 ( .A1(n564), .A2(n511), .ZN(n531) );
  NOR2_X1 U606 ( .A1(n509), .A2(n531), .ZN(n512) );
  XNOR2_X1 U607 ( .A(KEYINPUT28), .B(n512), .ZN(n513) );
  INV_X1 U608 ( .A(n534), .ZN(n584) );
  NAND2_X1 U609 ( .A1(n513), .A2(n584), .ZN(n526) );
  NAND2_X1 U610 ( .A1(n514), .A2(n679), .ZN(n515) );
  XNOR2_X2 U611 ( .A(n515), .B(KEYINPUT19), .ZN(n555) );
  INV_X1 U612 ( .A(n555), .ZN(n516) );
  NOR2_X1 U613 ( .A1(n526), .A2(n516), .ZN(n653) );
  INV_X1 U614 ( .A(n524), .ZN(n517) );
  NAND2_X1 U615 ( .A1(n525), .A2(n517), .ZN(n657) );
  INV_X1 U616 ( .A(n525), .ZN(n518) );
  NAND2_X1 U617 ( .A1(n524), .A2(n518), .ZN(n523) );
  NAND2_X1 U618 ( .A1(n657), .A2(n523), .ZN(n684) );
  NAND2_X1 U619 ( .A1(n653), .A2(n684), .ZN(n536) );
  NAND2_X1 U620 ( .A1(KEYINPUT47), .A2(n536), .ZN(n519) );
  NAND2_X1 U621 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U622 ( .A(KEYINPUT38), .B(n545), .ZN(n680) );
  NAND2_X1 U623 ( .A1(n507), .A2(n680), .ZN(n522) );
  NOR2_X1 U624 ( .A1(n525), .A2(n524), .ZN(n559) );
  INV_X1 U625 ( .A(n559), .ZN(n682) );
  XNOR2_X1 U626 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(n527), .ZN(n746) );
  NAND2_X1 U628 ( .A1(n744), .A2(n746), .ZN(n529) );
  XOR2_X1 U629 ( .A(KEYINPUT36), .B(n533), .Z(n535) );
  NOR2_X1 U630 ( .A1(KEYINPUT47), .A2(n536), .ZN(n537) );
  XNOR2_X1 U631 ( .A(n537), .B(KEYINPUT77), .ZN(n538) );
  INV_X1 U632 ( .A(n657), .ZN(n647) );
  AND2_X1 U633 ( .A1(n541), .A2(n647), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n542), .B(KEYINPUT108), .ZN(n745) );
  XOR2_X1 U635 ( .A(n349), .B(KEYINPUT104), .Z(n543) );
  NAND2_X1 U636 ( .A1(n543), .A2(n369), .ZN(n544) );
  XNOR2_X1 U637 ( .A(n544), .B(KEYINPUT43), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n546), .A2(n545), .ZN(n664) );
  INV_X1 U639 ( .A(n664), .ZN(n547) );
  OR2_X1 U640 ( .A1(n745), .A2(n547), .ZN(n548) );
  NOR2_X1 U641 ( .A1(G898), .A2(n736), .ZN(n728) );
  INV_X1 U642 ( .A(n550), .ZN(n551) );
  NAND2_X1 U643 ( .A1(n728), .A2(n551), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X2 U645 ( .A(n557), .B(n556), .ZN(n590) );
  INV_X1 U646 ( .A(n670), .ZN(n558) );
  AND2_X1 U647 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n590), .A2(n560), .ZN(n562) );
  AND2_X1 U649 ( .A1(n564), .A2(n509), .ZN(n563) );
  XNOR2_X1 U650 ( .A(n564), .B(KEYINPUT100), .ZN(n669) );
  NAND2_X1 U651 ( .A1(n669), .A2(n665), .ZN(n566) );
  XNOR2_X1 U652 ( .A(KEYINPUT101), .B(n566), .ZN(n567) );
  INV_X1 U653 ( .A(KEYINPUT32), .ZN(n568) );
  INV_X1 U654 ( .A(n743), .ZN(n569) );
  INV_X1 U655 ( .A(KEYINPUT65), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n577), .A2(n578), .ZN(n571) );
  XNOR2_X1 U657 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n572) );
  INV_X1 U658 ( .A(n590), .ZN(n586) );
  INV_X1 U659 ( .A(KEYINPUT34), .ZN(n574) );
  INV_X1 U660 ( .A(n577), .ZN(n580) );
  NOR2_X1 U661 ( .A1(n669), .A2(n581), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n636) );
  NAND2_X1 U663 ( .A1(n666), .A2(n584), .ZN(n585) );
  NOR2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n509), .A2(n587), .ZN(n642) );
  XOR2_X1 U666 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n592) );
  NAND2_X1 U667 ( .A1(n588), .A2(n484), .ZN(n589) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT93), .ZN(n675) );
  NAND2_X1 U669 ( .A1(n675), .A2(n590), .ZN(n591) );
  XNOR2_X1 U670 ( .A(n592), .B(n591), .ZN(n658) );
  NAND2_X1 U671 ( .A1(n642), .A2(n658), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n593), .A2(n684), .ZN(n594) );
  AND2_X1 U673 ( .A1(n636), .A2(n594), .ZN(n595) );
  XNOR2_X2 U674 ( .A(n596), .B(KEYINPUT45), .ZN(n720) );
  NAND2_X1 U675 ( .A1(n735), .A2(n720), .ZN(n702) );
  INV_X1 U676 ( .A(n702), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n597), .A2(n601), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n598), .A2(KEYINPUT85), .ZN(n605) );
  OR2_X1 U679 ( .A1(KEYINPUT85), .A2(n599), .ZN(n600) );
  NOR2_X1 U680 ( .A1(n702), .A2(n600), .ZN(n603) );
  AND2_X1 U681 ( .A1(n601), .A2(KEYINPUT2), .ZN(n602) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U683 ( .A(KEYINPUT86), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n735), .A2(KEYINPUT2), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n607), .B(n606), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n608), .A2(n720), .ZN(n704) );
  INV_X1 U687 ( .A(n629), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n609), .A2(G478), .ZN(n612) );
  INV_X1 U689 ( .A(G952), .ZN(n613) );
  AND2_X1 U690 ( .A1(n613), .A2(G953), .ZN(n719) );
  NAND2_X1 U691 ( .A1(n609), .A2(G210), .ZN(n621) );
  XNOR2_X1 U692 ( .A(KEYINPUT55), .B(KEYINPUT87), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT54), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U695 ( .A1(n622), .A2(n719), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U697 ( .A(G122), .B(KEYINPUT127), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(G24) );
  NOR2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT59), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U702 ( .A1(n633), .A2(n719), .ZN(n635) );
  XNOR2_X1 U703 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n634) );
  XNOR2_X1 U704 ( .A(n635), .B(n634), .ZN(G60) );
  XNOR2_X1 U705 ( .A(G101), .B(KEYINPUT110), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(G3) );
  INV_X1 U707 ( .A(n652), .ZN(n655) );
  NOR2_X1 U708 ( .A1(n642), .A2(n655), .ZN(n639) );
  XNOR2_X1 U709 ( .A(G104), .B(KEYINPUT111), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n641) );
  XNOR2_X1 U712 ( .A(G107), .B(KEYINPUT27), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n644) );
  NOR2_X1 U714 ( .A1(n657), .A2(n642), .ZN(n643) );
  XOR2_X1 U715 ( .A(n644), .B(n643), .Z(G9) );
  XNOR2_X1 U716 ( .A(n645), .B(G110), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT113), .ZN(G12) );
  XOR2_X1 U718 ( .A(G128), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U719 ( .A1(n653), .A2(n647), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U721 ( .A(G143), .B(n650), .Z(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT114), .B(n651), .ZN(G45) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(G146), .ZN(G48) );
  NOR2_X1 U725 ( .A1(n658), .A2(n655), .ZN(n656) );
  XOR2_X1 U726 ( .A(n348), .B(n656), .Z(G15) );
  NOR2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n660) );
  XNOR2_X1 U728 ( .A(G116), .B(KEYINPUT115), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(G18) );
  INV_X1 U730 ( .A(n661), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(G125), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U733 ( .A(G140), .B(n664), .ZN(G42) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT50), .B(n667), .Z(n668) );
  NAND2_X1 U736 ( .A1(n668), .A2(n509), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT49), .B(n671), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(KEYINPUT116), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n697), .A2(n678), .ZN(n692) );
  NOR2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(n683), .Z(n688) );
  INV_X1 U747 ( .A(n684), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n698), .A2(n689), .ZN(n690) );
  XNOR2_X1 U751 ( .A(n690), .B(KEYINPUT118), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n693), .Z(n694) );
  NAND2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT119), .ZN(n700) );
  NOR2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n706) );
  INV_X1 U758 ( .A(KEYINPUT2), .ZN(n701) );
  NAND2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U761 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(KEYINPUT120), .B(n707), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n708), .A2(G953), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n709), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U765 ( .A1(n716), .A2(G469), .ZN(n714) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  XOR2_X1 U767 ( .A(n710), .B(KEYINPUT121), .Z(n711) );
  XNOR2_X1 U768 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n714), .B(n713), .ZN(n715) );
  NOR2_X1 U770 ( .A1(n719), .A2(n715), .ZN(G54) );
  NOR2_X1 U771 ( .A1(n719), .A2(n718), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n720), .A2(n736), .ZN(n724) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n730) );
  XOR2_X1 U777 ( .A(n726), .B(n725), .Z(n727) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n731) );
  XOR2_X1 U780 ( .A(KEYINPUT125), .B(n731), .Z(G69) );
  XNOR2_X1 U781 ( .A(n732), .B(KEYINPUT126), .ZN(n733) );
  XOR2_X1 U782 ( .A(n734), .B(n733), .Z(n738) );
  XOR2_X1 U783 ( .A(n738), .B(n735), .Z(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U785 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U789 ( .A(G119), .B(n743), .Z(G21) );
  XNOR2_X1 U790 ( .A(G131), .B(n744), .ZN(G33) );
  XOR2_X1 U791 ( .A(G134), .B(n745), .Z(G36) );
  XNOR2_X1 U792 ( .A(G137), .B(n746), .ZN(G39) );
endmodule

