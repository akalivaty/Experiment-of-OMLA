//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT65), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  INV_X1    g014(.A(G96), .ZN(G221));
  INV_X1    g015(.A(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g027(.A1(G218), .A2(G221), .A3(G219), .ZN(new_n453));
  NAND3_X1  g028(.A1(new_n437), .A2(new_n438), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n456), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(new_n463), .B2(new_n462), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n469), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(G160));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n467), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n470), .A2(new_n471), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT71), .B1(new_n491), .B2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n481), .A2(new_n493), .A3(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(G124), .B2(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n470), .B2(new_n471), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(KEYINPUT72), .B(new_n500), .C1(new_n470), .C2(new_n471), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n467), .C1(new_n470), .C2(new_n471), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n481), .A2(new_n508), .A3(G138), .A4(new_n467), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n516), .A2(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G62), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n524), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n516), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n519), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n515), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n536), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  AOI22_X1  g117(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n525), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G90), .Z(new_n546));
  OAI22_X1  g121(.A1(new_n516), .A2(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n525), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n513), .A2(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n552));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n513), .B2(new_n514), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n552), .A2(G81), .B1(new_n554), .B2(G43), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G860), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n516), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n554), .A2(new_n567), .A3(new_n570), .A4(G53), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n571), .B1(G91), .B2(new_n552), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  INV_X1    g148(.A(G78), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n537), .A2(new_n573), .B1(new_n574), .B2(new_n553), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n577), .B1(new_n574), .B2(new_n553), .C1(new_n537), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(G651), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n572), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  OAI21_X1  g156(.A(KEYINPUT80), .B1(new_n524), .B2(new_n531), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n552), .A2(G88), .B1(new_n554), .B2(G50), .ZN(new_n583));
  INV_X1    g158(.A(G62), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n530), .B1(new_n537), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n582), .A2(new_n588), .ZN(G303));
  NAND2_X1  g164(.A1(new_n552), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n591));
  OAI211_X1 g166(.A(G49), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n552), .A2(G86), .B1(new_n554), .B2(G48), .ZN(new_n594));
  OAI21_X1  g169(.A(G61), .B1(new_n519), .B2(new_n518), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n525), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n525), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n516), .A2(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(G171), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n522), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT82), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n611), .B(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n537), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G54), .B2(new_n554), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n613), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n609), .B1(G868), .B2(new_n622), .ZN(G284));
  OAI21_X1  g198(.A(new_n609), .B1(G868), .B2(new_n622), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  INV_X1    g200(.A(G299), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  XNOR2_X1  g202(.A(G280), .B(KEYINPUT83), .ZN(G297));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND4_X1  g205(.A1(new_n613), .A2(new_n617), .A3(new_n629), .A4(new_n621), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(new_n558), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(G868), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n495), .A2(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(new_n486), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT84), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(G2096), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n643), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(G1341), .B(G1348), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT88), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT87), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n655), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT89), .Z(G401));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT90), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT17), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n676), .A2(KEYINPUT18), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n680), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT92), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n685), .B(new_n687), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n695), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n696), .A2(KEYINPUT20), .A3(new_n695), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n697), .B1(new_n695), .B2(new_n693), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G4), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n622), .B2(new_n711), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(G1348), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(G20), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT23), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G299), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1956), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(G1348), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n711), .A2(G19), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n633), .B2(new_n711), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1341), .Z(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT29), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n727), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G26), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n495), .A2(G128), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n737));
  INV_X1    g312(.A(G116), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G2105), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n640), .B2(G140), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2067), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n723), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G160), .A2(G29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G34), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n733), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n640), .A2(G139), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT25), .Z(new_n755));
  AOI22_X1  g330(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n755), .C1(new_n467), .C2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G33), .B(new_n757), .S(G29), .Z(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  NOR2_X1   g335(.A1(G171), .A2(new_n711), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G5), .B2(new_n711), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n727), .A2(G27), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G164), .B2(new_n727), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT100), .B(G2078), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n711), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n711), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n762), .A2(new_n760), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n724), .B1(new_n773), .B2(G28), .ZN(new_n775));
  AND2_X1   g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NOR2_X1   g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n642), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n727), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n771), .A2(new_n772), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n763), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n751), .A2(G2084), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n724), .A2(G32), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND3_X1  g361(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G141), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n787), .C1(new_n486), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G129), .B2(new_n495), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(new_n724), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT27), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1996), .ZN(new_n793));
  AND4_X1   g368(.A1(new_n752), .A2(new_n782), .A3(new_n783), .A4(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n720), .B(new_n744), .C1(new_n794), .C2(KEYINPUT101), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n711), .A2(G24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n605), .B2(new_n711), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1986), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n733), .A2(G25), .ZN(new_n799));
  INV_X1    g374(.A(G131), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n467), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n486), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G119), .B2(new_n495), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT95), .Z(new_n805));
  AOI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n727), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  AOI21_X1  g382(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n711), .A2(G6), .ZN(new_n809));
  INV_X1    g384(.A(G305), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n711), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G23), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  NOR3_X1   g391(.A1(new_n519), .A2(new_n518), .A3(G74), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n592), .B1(new_n817), .B2(new_n525), .ZN(new_n818));
  INV_X1    g393(.A(G87), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n522), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT98), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n590), .A2(new_n822), .A3(new_n591), .A4(new_n592), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n816), .B1(new_n824), .B2(new_n711), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n711), .A2(G22), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G166), .B2(new_n711), .ZN(new_n830));
  INV_X1    g405(.A(G1971), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n814), .A2(new_n827), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  OAI221_X1 g408(.A(new_n808), .B1(new_n806), .B2(new_n807), .C1(new_n833), .C2(KEYINPUT34), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(KEYINPUT34), .B2(new_n833), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  OR2_X1    g411(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n795), .A2(new_n836), .A3(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  AOI22_X1  g414(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n525), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n516), .A2(new_n842), .B1(new_n522), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n622), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT102), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  INV_X1    g425(.A(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n551), .A2(new_n557), .A3(new_n845), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT103), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n559), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(G160), .B(new_n642), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n486), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G130), .B2(new_n495), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n645), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n804), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n741), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n790), .B(new_n511), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n741), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n871), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n757), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT104), .Z(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n873), .B2(new_n876), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n862), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(new_n881), .A3(new_n886), .A4(new_n880), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g465(.A(KEYINPUT111), .B1(new_n851), .B2(new_n607), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n613), .A2(new_n617), .A3(new_n621), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G299), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n626), .A2(new_n613), .A3(new_n617), .A4(new_n621), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n895), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n852), .A2(new_n631), .A3(new_n853), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n631), .B1(new_n852), .B2(new_n853), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI211_X1 g481(.A(KEYINPUT108), .B(new_n899), .C1(new_n893), .C2(new_n895), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n898), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT42), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n824), .B(new_n605), .ZN(new_n916));
  XNOR2_X1  g491(.A(G166), .B(G305), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT109), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT110), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G868), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n912), .B2(new_n915), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n891), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n925), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(KEYINPUT111), .A3(G868), .A4(new_n923), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n926), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(G295));
  AND2_X1   g507(.A1(new_n926), .A2(new_n928), .ZN(G331));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n935));
  NAND2_X1  g510(.A1(G301), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n852), .B2(new_n853), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G286), .B1(G171), .B2(KEYINPUT113), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n852), .A2(new_n853), .A3(new_n936), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n902), .A2(new_n908), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n898), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n922), .ZN(new_n950));
  INV_X1    g525(.A(new_n922), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n898), .A2(new_n894), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n898), .B2(new_n899), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n941), .B2(new_n944), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n948), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n950), .A2(new_n955), .A3(new_n888), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n949), .B2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n945), .B2(new_n948), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n951), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n945), .A2(new_n948), .A3(new_n959), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n958), .B(new_n888), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n934), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n888), .B(new_n950), .C1(new_n961), .C2(new_n962), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n955), .A2(new_n888), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n965), .A2(KEYINPUT43), .B1(new_n966), .B2(new_n958), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n934), .ZN(G397));
  AOI21_X1  g543(.A(G1384), .B1(new_n505), .B2(new_n510), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G125), .ZN(new_n972));
  OR2_X1    g547(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n973));
  NAND2_X1  g548(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n473), .ZN(new_n976));
  OAI21_X1  g551(.A(G2105), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n483), .A2(G40), .A3(new_n977), .A4(new_n468), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n741), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n982), .B2(new_n790), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n980), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT46), .B1(new_n980), .B2(G1996), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n980), .A2(new_n982), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n988), .A2(KEYINPUT116), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(KEYINPUT116), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n790), .B(G1996), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n989), .B(new_n990), .C1(new_n980), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n807), .ZN(new_n993));
  OR3_X1    g568(.A1(new_n992), .A2(new_n805), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n874), .A2(new_n981), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n980), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n804), .B(new_n807), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n992), .B1(new_n979), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  AOI211_X1 g575(.A(new_n987), .B(new_n996), .C1(new_n998), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n511), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n978), .B1(new_n969), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n760), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT124), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n511), .B2(new_n1003), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n970), .A2(new_n1003), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n505), .B2(new_n510), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1011), .A2(new_n978), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G2078), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1004), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1013), .A2(new_n978), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1010), .A4(new_n1015), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT53), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1009), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT125), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT125), .B(new_n1009), .C1(new_n1016), .C2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n475), .A2(G40), .A3(new_n483), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n969), .B2(new_n970), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1017), .B(G1384), .C1(new_n505), .C2(new_n510), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1028), .A2(G2078), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(KEYINPUT53), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G301), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1028), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n969), .A2(KEYINPUT45), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(KEYINPUT53), .A3(new_n1015), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1009), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(new_n1031), .A3(G171), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1002), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G171), .B1(new_n1037), .B2(new_n1031), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT54), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1031), .A2(G171), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1041), .B1(new_n1026), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G8), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1027), .B2(new_n969), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n594), .A2(new_n598), .A3(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(G48), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n1048));
  INV_X1    g623(.A(G86), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n522), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(G1981), .B1(new_n1050), .B2(new_n597), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1051), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1045), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1045), .A2(new_n1054), .A3(KEYINPUT118), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n823), .A3(G1976), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1045), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1045), .B2(new_n1061), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n582), .A2(new_n588), .A3(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n831), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1005), .A2(new_n1007), .A3(new_n731), .ZN(new_n1074));
  AOI221_X4 g649(.A(new_n1044), .B1(new_n1071), .B2(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1006), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1004), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n969), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n731), .A3(new_n1080), .A4(new_n1027), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1076), .B1(new_n1082), .B2(G8), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1068), .A2(new_n1075), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G286), .A2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1013), .A2(new_n978), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n770), .B1(new_n1088), .B2(new_n1011), .ZN(new_n1089));
  INV_X1    g664(.A(G2084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1005), .A2(new_n1007), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1087), .B1(new_n1092), .B2(G8), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1005), .A2(new_n1007), .A3(new_n1090), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1966), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1091), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(G168), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1086), .A2(new_n1044), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1085), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1084), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1043), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n1105));
  XNOR2_X1  g680(.A(G299), .B(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1956), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1080), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1027), .B1(new_n969), .B2(new_n1006), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n971), .A2(new_n1027), .A3(new_n1035), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1008), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1027), .A2(new_n969), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G2067), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1119), .A3(new_n622), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n626), .A2(new_n1105), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1110), .A2(new_n1112), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1120), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1121), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1115), .A2(new_n892), .A3(new_n1118), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1348), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n622), .B1(new_n1130), .B2(new_n1117), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1119), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n892), .A2(KEYINPUT60), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1132), .A2(KEYINPUT60), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n971), .A2(new_n1137), .A3(new_n1027), .A4(new_n1035), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  AOI22_X1  g714(.A1(new_n1138), .A2(KEYINPUT121), .B1(new_n1116), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1034), .A2(new_n1141), .A3(new_n1137), .A4(new_n1035), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1143), .B2(new_n633), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT59), .B(new_n558), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1135), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1147), .C2(new_n1124), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n978), .B1(new_n1004), .B2(new_n1077), .ZN(new_n1150));
  AOI21_X1  g725(.A(G1956), .B1(new_n1150), .B2(new_n1080), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1111), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1028), .A2(new_n1029), .A3(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT122), .B(new_n1149), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1154), .B(new_n1155), .C1(new_n1156), .C2(new_n1113), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1148), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1128), .B1(new_n1146), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1039), .A2(new_n1104), .A3(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1044), .B(G286), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1084), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(KEYINPUT63), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1076), .B1(new_n1166), .B2(G8), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1162), .A2(new_n1163), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1075), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G288), .A2(G1976), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1060), .A2(new_n1171), .B1(new_n1046), .B2(new_n810), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1045), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1170), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1169), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1160), .A2(KEYINPUT126), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT126), .B1(new_n1160), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1033), .A2(new_n1180), .A3(new_n1084), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1101), .A2(KEYINPUT62), .A3(new_n1102), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1178), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n605), .B(G1986), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n998), .B1(new_n980), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1001), .B1(new_n1184), .B2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g762(.A1(new_n688), .A2(G319), .A3(new_n670), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1189), .A2(KEYINPUT127), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G229), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n889), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1193), .A2(new_n967), .ZN(G308));
  OR2_X1    g768(.A1(new_n1193), .A2(new_n967), .ZN(G225));
endmodule


