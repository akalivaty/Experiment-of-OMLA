//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT64), .B(G244), .Z(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND2_X1  g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G1), .A3(G13), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT66), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT66), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n244), .A2(new_n247), .A3(G1), .A4(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G222), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT65), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT65), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n250), .A2(new_n255), .A3(G222), .A4(new_n251), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n263), .A2(G223), .B1(G77), .B2(new_n262), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n249), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(new_n245), .A3(G274), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n245), .A2(new_n266), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n214), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n206), .A2(G33), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR3_X1   g0082(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n276), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT68), .B1(new_n206), .B2(G1), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n205), .A3(G20), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n276), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(new_n296), .B1(new_n292), .B2(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n265), .B2(new_n271), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n274), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n272), .A2(G190), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n272), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n298), .B(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT72), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n298), .B(KEYINPUT70), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT9), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT71), .B1(new_n310), .B2(KEYINPUT9), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n307), .A2(new_n315), .A3(new_n308), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n313), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n302), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n295), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT12), .ZN(new_n325));
  INV_X1    g0125(.A(new_n291), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G68), .A3(new_n296), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n284), .A2(new_n292), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n278), .A2(new_n218), .B1(new_n206), .B2(G68), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n276), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT11), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n331), .B(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n259), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n250), .A2(KEYINPUT73), .A3(G232), .A4(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n250), .A2(G226), .A3(new_n251), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n249), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G238), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n268), .B1(new_n269), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n341), .B2(new_n342), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(G190), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n331), .B(KEYINPUT11), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n334), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n348), .A2(new_n357), .A3(new_n351), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n349), .A2(KEYINPUT74), .A3(new_n350), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n360), .B2(G200), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(G169), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n358), .A2(new_n364), .A3(G169), .A4(new_n359), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n348), .A2(G179), .A3(new_n351), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n334), .A2(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(new_n323), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n284), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n258), .A2(KEYINPUT76), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G33), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT3), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n258), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n376), .B(new_n206), .C1(new_n380), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT3), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n260), .ZN(new_n388));
  NAND2_X1  g0188(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G33), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(G20), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n376), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT16), .B(new_n375), .C1(new_n385), .C2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n376), .A2(G20), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT3), .B1(new_n377), .B2(new_n379), .ZN(new_n396));
  AOI21_X1  g0196(.A(G33), .B1(new_n388), .B2(new_n389), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n376), .B1(new_n250), .B2(G20), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n323), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n394), .B1(new_n400), .B2(new_n374), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(new_n401), .A3(new_n276), .ZN(new_n402));
  INV_X1    g0202(.A(new_n279), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n326), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n296), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n294), .B2(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n270), .B2(G1698), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n386), .A2(new_n410), .A3(new_n390), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n342), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n268), .B1(new_n269), .B2(new_n229), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n299), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n249), .B1(new_n411), .B2(new_n412), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n418), .A2(new_n273), .A3(new_n415), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n408), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n408), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G190), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(KEYINPUT79), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(KEYINPUT79), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n414), .A2(new_n416), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n304), .B1(new_n418), .B2(new_n415), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n402), .A2(new_n433), .A3(new_n407), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n402), .A2(new_n433), .A3(KEYINPUT17), .A4(new_n407), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n291), .A2(new_n218), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n296), .B1(new_n218), .B2(new_n295), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n284), .A2(new_n279), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n443), .A2(new_n278), .B1(new_n206), .B2(new_n218), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n276), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT69), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n263), .A2(G238), .B1(G107), .B2(new_n262), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n229), .B2(new_n252), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n342), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n269), .A2(new_n217), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n245), .A2(G274), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n266), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n448), .B(new_n457), .C1(new_n426), .C2(new_n456), .ZN(new_n458));
  INV_X1    g0258(.A(new_n446), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n456), .B2(new_n299), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G179), .B2(new_n456), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n322), .A2(new_n369), .A3(new_n439), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n294), .A2(G97), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n296), .B1(G1), .B2(new_n258), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G97), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n469), .A2(KEYINPUT6), .ZN(new_n470));
  INV_X1    g0270(.A(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(KEYINPUT80), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G107), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n470), .A2(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g0278(.A(G20), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n284), .A2(new_n218), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(KEYINPUT81), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n472), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n473), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n206), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n487), .B2(new_n480), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n398), .A2(new_n399), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G107), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n482), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n468), .B1(new_n491), .B2(new_n276), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n494), .A2(new_n245), .A3(G274), .A4(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n245), .ZN(new_n501));
  INV_X1    g0301(.A(G257), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G244), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(G1698), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n386), .A2(new_n390), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT4), .A2(G244), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n259), .A2(new_n261), .A3(new_n509), .A4(new_n251), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n259), .A2(new_n261), .A3(G250), .A4(G1698), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n503), .B1(new_n514), .B2(new_n342), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G169), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n497), .B(new_n518), .C1(new_n501), .C2(new_n502), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n249), .B1(new_n508), .B2(new_n513), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n273), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n493), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n491), .A2(new_n276), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(G190), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n525), .A2(new_n467), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT25), .ZN(new_n530));
  AOI211_X1 g0330(.A(G107), .B(new_n294), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G107), .B2(new_n466), .ZN(new_n535));
  NOR2_X1   g0335(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n471), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT84), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n377), .A2(new_n379), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n206), .A3(G116), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n541), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n386), .A2(new_n390), .A3(new_n206), .A4(G87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT22), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n206), .A3(G87), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n262), .A2(KEYINPUT83), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  INV_X1    g0353(.A(G87), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n554), .A2(KEYINPUT22), .A3(G20), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n250), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n537), .B1(new_n547), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n541), .A2(new_n544), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT84), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n541), .A2(new_n544), .A3(new_n542), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n549), .A2(new_n557), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n536), .A4(new_n538), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n276), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n535), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G250), .A2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n502), .B2(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n386), .A2(new_n570), .A3(new_n390), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n543), .A2(G294), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n500), .A2(new_n245), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n573), .A2(new_n342), .B1(G264), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n497), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(G190), .A3(new_n497), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n524), .B(new_n528), .C1(new_n568), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n576), .A2(G179), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n575), .B2(new_n497), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n567), .B1(new_n559), .B2(new_n565), .ZN(new_n584));
  INV_X1    g0384(.A(new_n535), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n512), .B(new_n206), .C1(G33), .C2(new_n469), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n276), .C1(new_n206), .C2(G116), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT20), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n296), .B(G116), .C1(G1), .C2(new_n258), .ZN(new_n591));
  INV_X1    g0391(.A(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n295), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  MUX2_X1   g0395(.A(G257), .B(G264), .S(G1698), .Z(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n386), .A3(new_n390), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n262), .A2(G303), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n249), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n500), .A2(G270), .A3(new_n245), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n497), .ZN(new_n601));
  OAI21_X1  g0401(.A(G169), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n587), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(G200), .B1(new_n599), .B2(new_n601), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n599), .A2(new_n601), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n595), .B(new_n604), .C1(new_n605), .C2(new_n430), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n599), .A2(new_n273), .A3(new_n601), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n589), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n589), .A2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n593), .B(new_n591), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(new_n611), .A3(KEYINPUT21), .A4(G169), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n603), .A2(new_n606), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n386), .A2(new_n390), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n206), .A3(G68), .ZN(new_n616));
  NOR3_X1   g0416(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n206), .B2(new_n339), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G97), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n618), .A2(new_n619), .B1(new_n278), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n276), .ZN(new_n623));
  INV_X1    g0423(.A(new_n443), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n294), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n466), .A2(new_n624), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n205), .A2(G45), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n245), .A2(G250), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n453), .B2(new_n629), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n543), .A2(G116), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n386), .A2(new_n390), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n344), .A2(new_n251), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n504), .A2(G1698), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n631), .B1(new_n637), .B2(new_n342), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n273), .ZN(new_n639));
  INV_X1    g0439(.A(new_n638), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n299), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n628), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n567), .B1(new_n616), .B2(new_n621), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n465), .A2(new_n554), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n643), .A2(new_n625), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(G200), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(G190), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n586), .A2(new_n614), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n463), .A2(new_n580), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT87), .ZN(G372));
  NAND2_X1  g0452(.A1(new_n319), .A2(new_n321), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n361), .A2(new_n461), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n367), .A2(new_n368), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n438), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n656), .B2(new_n425), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n301), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n386), .A2(new_n390), .A3(new_n634), .A4(new_n635), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n249), .B1(new_n660), .B2(new_n632), .ZN(new_n661));
  OAI211_X1 g0461(.A(KEYINPUT88), .B(new_n299), .C1(new_n661), .C2(new_n631), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n638), .B2(G169), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT89), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(KEYINPUT89), .A3(new_n639), .A4(new_n662), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n628), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n648), .ZN(new_n671));
  INV_X1    g0471(.A(new_n628), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n665), .A2(new_n639), .A3(new_n662), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT89), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n672), .B1(new_n675), .B2(new_n667), .ZN(new_n676));
  INV_X1    g0476(.A(new_n648), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT90), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  INV_X1    g0480(.A(new_n524), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n603), .A2(new_n613), .A3(new_n612), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n568), .B2(new_n583), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n580), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  AND4_X1   g0486(.A1(new_n493), .A2(new_n523), .A3(new_n648), .A4(new_n642), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n669), .B1(new_n687), .B2(new_n680), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n682), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n659), .B1(new_n463), .B2(new_n691), .ZN(G369));
  NOR3_X1   g0492(.A1(new_n584), .A2(new_n579), .A3(new_n585), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n693), .B1(new_n568), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n586), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n611), .A2(new_n699), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  MUX2_X1   g0508(.A(new_n614), .B(new_n683), .S(new_n708), .Z(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n700), .A2(new_n701), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n683), .A2(new_n703), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n705), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(G41), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n209), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n617), .A2(new_n592), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n212), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT94), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n670), .B1(new_n669), .B2(new_n648), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n676), .A2(KEYINPUT90), .A3(new_n677), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n681), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT26), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n676), .B1(new_n687), .B2(new_n680), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT95), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n685), .A2(new_n679), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n728), .A2(new_n732), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n688), .B1(new_n685), .B2(new_n679), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n699), .B1(new_n738), .B2(new_n682), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(KEYINPUT29), .B2(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n586), .A2(new_n614), .A3(new_n649), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n517), .A2(new_n519), .ZN(new_n742));
  INV_X1    g0542(.A(new_n521), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n744), .A2(G179), .B1(G169), .B2(new_n515), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n528), .B1(new_n745), .B2(new_n492), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n693), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n747), .A3(new_n703), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n515), .A2(new_n607), .A3(new_n575), .A4(new_n638), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n638), .A2(new_n575), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n515), .A4(new_n607), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n742), .A2(new_n743), .B1(new_n575), .B2(new_n497), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n640), .A2(new_n605), .A3(new_n273), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n699), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n751), .A2(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n703), .A2(new_n761), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(G330), .B1(new_n749), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n740), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n727), .B1(new_n768), .B2(G1), .ZN(G364));
  INV_X1    g0569(.A(new_n720), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n206), .A2(G13), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n205), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n710), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G330), .B2(new_n709), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n209), .A2(new_n250), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n778), .B1(G116), .B2(new_n209), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n239), .A2(new_n495), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n633), .A2(new_n209), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n495), .B2(new_n213), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n214), .B1(G20), .B2(new_n299), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n774), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(G20), .A2(G179), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n429), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G322), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n426), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n206), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n792), .A2(new_n426), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(G311), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n304), .A2(G179), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(G20), .A3(new_n426), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(G20), .A3(G190), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n206), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n250), .B(new_n808), .C1(G329), .C2(new_n809), .ZN(new_n810));
  OR3_X1    g0610(.A1(new_n791), .A2(new_n304), .A3(KEYINPUT96), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT96), .B1(new_n791), .B2(new_n304), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n429), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n811), .A2(new_n426), .A3(new_n812), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n814), .A2(G326), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n802), .A2(new_n810), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n809), .A2(G159), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n794), .A2(new_n370), .B1(KEYINPUT32), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G77), .B2(new_n801), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n250), .B1(new_n806), .B2(new_n554), .ZN(new_n823));
  INV_X1    g0623(.A(new_n804), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(G107), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n798), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G97), .B1(new_n820), .B2(KEYINPUT32), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n822), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n813), .A2(new_n292), .B1(new_n815), .B2(new_n323), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n790), .B1(new_n830), .B2(new_n787), .ZN(new_n831));
  INV_X1    g0631(.A(new_n786), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n709), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n776), .A2(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n690), .A2(new_n703), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n458), .B1(new_n459), .B2(new_n703), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n461), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n461), .A2(new_n699), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n739), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(new_n767), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n774), .B1(new_n844), .B2(new_n767), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n774), .ZN(new_n848));
  INV_X1    g0648(.A(new_n787), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n793), .A2(G143), .B1(G159), .B2(new_n801), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n851), .B2(new_n813), .C1(new_n285), .C2(new_n815), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT34), .ZN(new_n853));
  INV_X1    g0653(.A(new_n809), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(new_n292), .B2(new_n806), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G68), .B2(new_n824), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n633), .B1(new_n826), .B2(G58), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n814), .A2(G303), .B1(G283), .B2(new_n816), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n250), .B1(new_n809), .B2(G311), .ZN(new_n861));
  INV_X1    g0661(.A(new_n806), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n862), .A2(G107), .B1(new_n824), .B2(G87), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n798), .A2(new_n469), .B1(new_n800), .B2(new_n592), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n793), .B2(G294), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n860), .A2(new_n861), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n849), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n787), .A2(new_n784), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n848), .B(new_n867), .C1(new_n218), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n842), .B2(new_n785), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT97), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n847), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n477), .A2(new_n478), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(G116), .A3(new_n215), .A4(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT36), .Z(new_n879));
  OR3_X1    g0679(.A1(new_n212), .A2(new_n218), .A3(new_n371), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n292), .A2(G68), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n205), .B(G13), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n323), .B1(new_n391), .B2(new_n376), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT7), .B1(new_n615), .B2(G20), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n374), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n567), .B1(new_n886), .B2(KEYINPUT16), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n375), .B1(new_n385), .B2(new_n392), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n394), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n406), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT98), .B1(new_n890), .B2(new_n697), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n393), .A2(new_n276), .ZN(new_n892));
  INV_X1    g0692(.A(new_n394), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n884), .A2(new_n885), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n375), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n407), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT98), .ZN(new_n897));
  INV_X1    g0697(.A(new_n697), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n420), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n891), .A2(new_n434), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT99), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n434), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n417), .A2(new_n419), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n402), .A2(new_n407), .B1(new_n906), .B2(new_n697), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n393), .A2(new_n401), .A3(new_n276), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(new_n406), .B1(new_n420), .B2(new_n898), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(KEYINPUT99), .A3(new_n904), .A4(new_n434), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n393), .B(new_n276), .C1(new_n886), .C2(new_n893), .ZN(new_n914));
  AOI211_X1 g0714(.A(KEYINPUT98), .B(new_n697), .C1(new_n914), .C2(new_n407), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n425), .A2(new_n438), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n901), .A2(KEYINPUT37), .B1(new_n908), .B2(new_n911), .ZN(new_n919));
  AOI211_X1 g0719(.A(KEYINPUT18), .B(new_n906), .C1(new_n402), .C2(new_n407), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n423), .B1(new_n408), .B2(new_n420), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n436), .A2(new_n437), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n923), .B1(new_n899), .B2(new_n891), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n919), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT39), .B1(new_n918), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n915), .A2(new_n916), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n900), .A2(new_n434), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n904), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n908), .A2(new_n911), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT38), .B(new_n917), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT100), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n434), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n402), .A2(new_n433), .A3(KEYINPUT100), .A4(new_n407), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n910), .A3(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n908), .A2(new_n911), .B1(new_n936), .B2(KEYINPUT37), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n408), .A2(new_n898), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n922), .B2(new_n923), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n925), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n927), .B(KEYINPUT101), .C1(KEYINPUT39), .C2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n655), .A2(new_n699), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT101), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n932), .A2(new_n940), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n425), .A2(new_n697), .ZN(new_n948));
  INV_X1    g0748(.A(new_n361), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n368), .A2(new_n699), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n655), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n368), .B(new_n699), .C1(new_n367), .C2(new_n361), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n699), .B(new_n840), .C1(new_n738), .C2(new_n682), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n953), .B1(new_n926), .B2(new_n918), .C1(new_n954), .C2(new_n838), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n948), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT29), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n463), .B1(new_n835), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n737), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT102), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT102), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n737), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n658), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n957), .B(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(G330), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT103), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n759), .A2(new_n967), .A3(new_n764), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT103), .B1(new_n763), .B2(new_n765), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n968), .A2(new_n969), .B1(new_n760), .B2(new_n761), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n748), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n463), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT104), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n840), .B1(new_n970), .B2(new_n748), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n912), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n408), .B(new_n898), .C1(new_n425), .C2(new_n438), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT38), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n953), .B(new_n975), .C1(new_n926), .C2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n975), .A2(new_n953), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n925), .B1(new_n919), .B2(new_n924), .ZN(new_n982));
  AOI21_X1  g0782(.A(KEYINPUT40), .B1(new_n982), .B2(new_n932), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n980), .A2(KEYINPUT40), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n966), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n974), .B2(new_n985), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n965), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n205), .B2(new_n771), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n965), .A2(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n883), .B1(new_n989), .B2(new_n990), .ZN(G367));
  OAI221_X1 g0791(.A(new_n788), .B1(new_n209), .B2(new_n443), .C1(new_n235), .C2(new_n781), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n992), .A2(new_n774), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n826), .A2(G68), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n794), .B2(new_n285), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G50), .B2(new_n801), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n804), .A2(new_n218), .B1(new_n806), .B2(new_n370), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n262), .B(new_n997), .C1(G137), .C2(new_n809), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n814), .A2(G143), .B1(G159), .B2(new_n816), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n806), .A2(new_n592), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(KEYINPUT46), .B1(new_n805), .B2(new_n800), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT46), .B2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n804), .A2(new_n469), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1004), .B(new_n615), .C1(G317), .C2(new_n809), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n793), .A2(G303), .B1(G107), .B2(new_n826), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G311), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n813), .A2(new_n1008), .B1(new_n815), .B2(new_n796), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n645), .A2(new_n703), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n679), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n669), .A2(new_n1013), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n993), .B1(new_n849), .B2(new_n1012), .C1(new_n1017), .C2(new_n832), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT108), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n681), .A2(new_n699), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n524), .B(new_n528), .C1(new_n492), .C2(new_n703), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n717), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT45), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n717), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n717), .B2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT106), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n713), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n712), .B(KEYINPUT106), .C1(new_n1024), .C2(new_n1029), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n706), .B(new_n716), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(new_n710), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n768), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n768), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n720), .B(KEYINPUT41), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n773), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n706), .A2(new_n716), .A3(new_n1022), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(KEYINPUT42), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n524), .B1(new_n1021), .B2(new_n586), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n703), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1041), .A2(KEYINPUT42), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT43), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1016), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1017), .A2(KEYINPUT43), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1045), .A2(new_n1048), .A3(new_n1016), .A4(new_n1046), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n712), .A2(new_n1022), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1019), .B1(new_n1040), .B2(new_n1055), .ZN(G387));
  OAI22_X1  g0856(.A1(new_n777), .A2(new_n722), .B1(G107), .B2(new_n209), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n232), .A2(new_n495), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n279), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n721), .C1(G68), .C2(G77), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n781), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n774), .B1(new_n789), .B2(new_n1063), .C1(new_n706), .C2(new_n832), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n793), .A2(G317), .B1(G303), .B2(new_n801), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n1008), .B2(new_n815), .C1(new_n795), .C2(new_n813), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n826), .A2(G283), .B1(new_n862), .B2(G294), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT49), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT109), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n824), .A2(G116), .B1(new_n809), .B2(G326), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n633), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n814), .A2(G159), .B1(new_n403), .B2(new_n816), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n806), .A2(new_n218), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1078), .B(new_n1004), .C1(G150), .C2(new_n809), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n798), .A2(new_n443), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(new_n633), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n793), .A2(G50), .B1(G68), .B2(new_n801), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1064), .B1(new_n1084), .B2(new_n787), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1035), .B2(new_n773), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1036), .A2(new_n770), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n768), .A2(new_n1035), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(G393));
  NAND2_X1  g0889(.A1(new_n713), .A2(KEYINPUT110), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT110), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n712), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(new_n1024), .C2(new_n1029), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n1091), .A3(new_n712), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n773), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n788), .B1(new_n469), .B2(new_n209), .C1(new_n242), .C2(new_n781), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n774), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n862), .A2(G283), .B1(G322), .B2(new_n809), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n262), .C1(new_n471), .C2(new_n804), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT111), .Z(new_n1102));
  AOI22_X1  g0902(.A1(new_n826), .A2(G116), .B1(new_n801), .B2(G294), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n807), .C2(new_n815), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n814), .A2(G317), .B1(new_n793), .B2(G311), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT52), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n814), .A2(G150), .B1(new_n793), .B2(G159), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n798), .A2(new_n218), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n633), .B(new_n1109), .C1(new_n403), .C2(new_n801), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n804), .A2(new_n554), .B1(new_n806), .B2(new_n323), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G143), .B2(new_n809), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(new_n292), .C2(new_n815), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1104), .A2(new_n1106), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1099), .B1(new_n1114), .B2(new_n787), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1022), .B2(new_n832), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1096), .B1(new_n768), .B2(new_n1035), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n770), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1097), .B(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(G390));
  NOR3_X1   g0919(.A1(new_n463), .A2(new_n972), .A3(new_n966), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n959), .A2(new_n737), .A3(new_n962), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n962), .B1(new_n959), .B2(new_n737), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n659), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n736), .A2(new_n703), .A3(new_n837), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1126), .A2(new_n839), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n953), .B1(G330), .B2(new_n975), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n767), .A2(new_n840), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n953), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n838), .B1(new_n739), .B2(new_n842), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n975), .A2(new_n953), .A3(G330), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1129), .B2(new_n953), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1134), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n943), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n953), .B1(new_n954), .B2(new_n838), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n942), .B2(new_n946), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n941), .A2(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1126), .A2(new_n839), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n953), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1139), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n953), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1140), .B1(new_n1132), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT101), .B1(new_n941), .B2(KEYINPUT39), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n945), .B1(new_n982), .B2(new_n932), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n946), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1129), .A2(new_n953), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1147), .B1(new_n1126), .B2(new_n839), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1153), .C1(new_n1154), .C2(new_n1143), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1146), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1138), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1125), .A2(new_n1146), .A3(new_n1155), .A4(new_n1137), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n770), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n784), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n868), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n774), .B1(new_n403), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n800), .A2(new_n469), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1109), .B(new_n1164), .C1(new_n793), .C2(G116), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n814), .A2(G283), .B1(G107), .B2(new_n816), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n250), .B1(new_n862), .B2(G87), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n824), .A2(G68), .B1(new_n809), .B2(G294), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n285), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT53), .B1(new_n806), .B2(new_n285), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n794), .B2(new_n855), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G159), .C2(new_n826), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT54), .B(G143), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n815), .A2(new_n851), .B1(new_n800), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT112), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n814), .A2(G128), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n804), .A2(new_n292), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n262), .B(new_n1178), .C1(G125), .C2(new_n809), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1175), .A2(KEYINPUT112), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1169), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1163), .B1(new_n1182), .B2(new_n787), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1160), .A2(new_n773), .B1(new_n1161), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1159), .A2(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(KEYINPUT117), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT116), .B1(new_n984), .B2(new_n966), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT116), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n981), .A2(new_n983), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT40), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n981), .B2(new_n941), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(G330), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n310), .A2(new_n697), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n322), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n322), .A2(new_n1196), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1194), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1199), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1197), .A3(new_n1193), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1187), .A2(new_n1192), .A3(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(KEYINPUT116), .C1(new_n984), .C2(new_n966), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1205), .A2(new_n956), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n956), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1186), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n957), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(new_n956), .A3(new_n1206), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(KEYINPUT117), .A3(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1127), .A2(new_n1130), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1125), .B1(new_n1156), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(new_n1158), .B2(new_n1125), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n720), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1209), .A2(new_n1213), .A3(new_n773), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n848), .B1(new_n292), .B2(new_n868), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n615), .A2(G41), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G33), .A2(G41), .ZN(new_n1226));
  OR3_X1    g1026(.A1(new_n1225), .A2(G50), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n804), .A2(new_n370), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1078), .B(new_n1228), .C1(G283), .C2(new_n809), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n793), .A2(G107), .B1(new_n624), .B2(new_n801), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1225), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n994), .B1(new_n813), .B2(new_n592), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT113), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G97), .C2(new_n816), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1227), .B1(new_n1234), .B2(KEYINPUT58), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT114), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n814), .A2(G125), .B1(G132), .B2(new_n816), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n806), .A2(new_n1174), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT115), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n826), .A2(G150), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n793), .A2(G128), .B1(G137), .B2(new_n801), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n809), .A2(G124), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1226), .C1(new_n373), .C2(new_n804), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1242), .B2(KEYINPUT59), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1234), .A2(KEYINPUT58), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1236), .A2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1224), .B1(new_n849), .B2(new_n1248), .C1(new_n1203), .C2(new_n785), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1223), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1222), .A2(new_n1251), .ZN(G375));
  INV_X1    g1052(.A(KEYINPUT119), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1137), .A2(new_n1253), .A3(new_n773), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT119), .B1(new_n1214), .B2(new_n772), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n774), .B1(G68), .B2(new_n1162), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n794), .A2(new_n851), .B1(new_n292), .B2(new_n798), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G150), .B2(new_n801), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n809), .A2(G128), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n373), .B2(new_n806), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n633), .B(new_n1228), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n815), .A2(new_n1174), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1258), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n813), .A2(new_n855), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT121), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1080), .B1(new_n793), .B2(G283), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n1269), .A2(KEYINPUT120), .B1(G294), .B2(new_n814), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(KEYINPUT120), .B2(new_n1269), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n854), .A2(new_n807), .B1(new_n469), .B2(new_n806), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n250), .B(new_n1272), .C1(G77), .C2(new_n824), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n471), .B2(new_n800), .C1(new_n592), .C2(new_n815), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1265), .A2(new_n1267), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1256), .B1(new_n1275), .B2(new_n787), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n953), .B2(new_n785), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1254), .A2(new_n1255), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1124), .A2(new_n1214), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1038), .B(KEYINPUT118), .Z(new_n1281));
  NAND3_X1  g1081(.A1(new_n1138), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(G381));
  NOR2_X1   g1083(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1097), .A2(new_n1116), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n872), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G396), .A2(new_n1287), .A3(G387), .A4(G393), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G378), .A2(new_n1288), .A3(G375), .A4(G381), .ZN(G407));
  AOI21_X1  g1089(.A(new_n1250), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1290));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n698), .A2(G213), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1293), .ZN(G409));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1222), .A2(G378), .A3(new_n1251), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1209), .A2(new_n1213), .A3(new_n1215), .A4(new_n1281), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1249), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1220), .B2(new_n773), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G378), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1292), .B1(new_n1296), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1214), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1303), .A2(new_n770), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1124), .A2(new_n1214), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1280), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1279), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n872), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(G384), .A3(new_n1279), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1292), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1308), .B2(new_n1279), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n872), .B(new_n1278), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1313), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1315), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1295), .B1(new_n1302), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT124), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1302), .A2(KEYINPUT63), .A3(new_n1318), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1321), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1300), .B1(new_n1290), .B2(G378), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(new_n1325), .A2(new_n1326), .A3(new_n1292), .A4(new_n1312), .ZN(new_n1327));
  XOR2_X1   g1127(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1302), .B2(new_n1318), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT124), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(new_n1286), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G390), .B(new_n1019), .C1(new_n1040), .C2(new_n1055), .ZN(new_n1333));
  XOR2_X1   g1133(.A(G393), .B(G396), .Z(new_n1334));
  AND3_X1   g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1334), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT125), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1339), .B(new_n1295), .C1(new_n1302), .C2(new_n1320), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1316), .A2(new_n1317), .A3(new_n1314), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1313), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1325), .B2(new_n1292), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT125), .B1(new_n1345), .B2(new_n1295), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1341), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1302), .A2(new_n1318), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1302), .B(new_n1318), .C1(KEYINPUT126), .C2(KEYINPUT62), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  AOI22_X1  g1153(.A1(new_n1331), .A2(new_n1337), .B1(new_n1347), .B2(new_n1353), .ZN(G405));
  OAI21_X1  g1154(.A(new_n1312), .B1(new_n1290), .B2(G378), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(G375), .A2(new_n1291), .A3(new_n1318), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1357), .A2(KEYINPUT127), .A3(new_n1296), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1355), .A2(new_n1356), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1358), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1337), .ZN(new_n1362));
  XNOR2_X1  g1162(.A(new_n1361), .B(new_n1362), .ZN(G402));
endmodule


