//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(KEYINPUT66), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT27), .B(G183gat), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n211), .A2(new_n212), .A3(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  AOI21_X1  g014(.A(G190gat), .B1(new_n215), .B2(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  OR3_X1    g016(.A1(new_n217), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT28), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n209), .B(new_n210), .C1(new_n213), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n221), .A2(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n222), .A2(new_n225), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n217), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n232), .A2(KEYINPUT24), .A3(new_n210), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n230), .A2(new_n233), .B1(KEYINPUT64), .B2(new_n221), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n222), .A2(new_n229), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n225), .A2(new_n227), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(KEYINPUT24), .A3(new_n210), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G120gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G134gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n249), .B2(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n247), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(KEYINPUT67), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n220), .A2(new_n240), .A3(new_n253), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G227gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT34), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n257), .A2(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G71gat), .ZN(new_n266));
  INV_X1    g065(.A(G99gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n260), .A3(new_n256), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT33), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n262), .A2(new_n263), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n271), .B(KEYINPUT32), .C1(new_n272), .C2(new_n270), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n277), .B1(new_n275), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n265), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n276), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n264), .A3(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G22gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G162gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G155gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G141gat), .B(G148gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n297));
  XNOR2_X1  g096(.A(G155gat), .B(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n295), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT76), .B(G155gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n303), .B2(new_n290), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n301), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT22), .ZN(new_n311));
  NAND2_X1  g110(.A1(G211gat), .A2(G218gat), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  OR2_X1    g114(.A1(G211gat), .A2(G218gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n312), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n315), .A3(new_n312), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n319), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n313), .B1(new_n321), .B2(new_n317), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n322), .A3(KEYINPUT71), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n318), .A2(new_n314), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n308), .B1(new_n327), .B2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n325), .ZN(new_n331));
  INV_X1    g130(.A(new_n296), .ZN(new_n332));
  INV_X1    g131(.A(new_n295), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n298), .A2(new_n299), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n304), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT77), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI211_X1 g137(.A(KEYINPUT3), .B(new_n332), .C1(new_n338), .C2(new_n305), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n331), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n340));
  INV_X1    g139(.A(G228gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(new_n259), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n308), .B(KEYINPUT81), .C1(new_n327), .C2(KEYINPUT3), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n330), .A2(new_n340), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n331), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n296), .C1(new_n306), .C2(new_n307), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n347), .B2(new_n326), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n332), .B1(new_n338), .B2(new_n305), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n320), .A2(new_n322), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n326), .C1(new_n350), .C2(new_n322), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n348), .A2(new_n353), .B1(new_n341), .B2(new_n259), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT31), .B(G50gat), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n344), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n344), .B2(new_n354), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n289), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n354), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n354), .A3(new_n356), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n288), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n202), .B1(new_n286), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n366), .B(KEYINPUT72), .Z(new_n367));
  NAND2_X1  g166(.A1(new_n241), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n241), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n220), .A2(new_n240), .A3(KEYINPUT73), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n345), .B(new_n368), .C1(new_n372), .C2(new_n367), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n367), .A2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n241), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  INV_X1    g175(.A(new_n367), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n331), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n378), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n383), .A2(KEYINPUT30), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n254), .B1(new_n308), .B2(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n347), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n349), .A2(new_n254), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n332), .B(new_n253), .C1(new_n338), .C2(new_n305), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n391), .A2(new_n392), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n308), .A2(new_n253), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(new_n392), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n394), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n349), .A2(new_n254), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n396), .B2(KEYINPUT4), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT5), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n402), .B1(new_n390), .B2(new_n347), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n398), .A2(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(G1gat), .B(G29gat), .Z(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n403), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n407), .A2(new_n408), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n389), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n281), .A2(new_n285), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n424), .A2(KEYINPUT85), .A3(new_n363), .A4(new_n359), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n365), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n286), .A2(new_n364), .A3(KEYINPUT35), .ZN(new_n428));
  INV_X1    g227(.A(new_n389), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n414), .B1(new_n409), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n416), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n422), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n431), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n253), .B1(new_n349), .B2(new_n346), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n339), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n441), .B(new_n402), .C1(new_n443), .C2(new_n406), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n415), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n447), .A3(new_n415), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n402), .B1(new_n443), .B2(new_n406), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(KEYINPUT39), .C1(new_n402), .C2(new_n401), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n440), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n444), .A2(new_n447), .A3(new_n415), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n444), .B2(new_n415), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n440), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n389), .B(new_n439), .C1(new_n452), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n364), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n385), .B1(new_n384), .B2(KEYINPUT37), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n373), .B2(new_n378), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT38), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n382), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n376), .A2(new_n377), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n464), .B1(new_n241), .B2(new_n374), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n460), .B1(new_n465), .B2(new_n345), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n331), .B(new_n368), .C1(new_n372), .C2(new_n367), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n459), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n434), .A2(new_n422), .A3(new_n462), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n457), .A2(new_n458), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n424), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n281), .A2(new_n285), .A3(KEYINPUT36), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n359), .A2(new_n363), .A3(KEYINPUT82), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT82), .B1(new_n359), .B2(new_n363), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n421), .A2(new_n422), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n429), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n437), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(G197gat), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT11), .B(G169gat), .Z(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT12), .Z(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(G43gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(G50gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(G43gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n496), .A2(G43gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(G50gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT15), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NOR2_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n512), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n492), .B1(new_n507), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT15), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT15), .B1(new_n504), .B2(new_n505), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR4_X1   g321(.A1(KEYINPUT88), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n515), .B2(new_n512), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n508), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT89), .A4(new_n503), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT90), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n508), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n503), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n529), .A2(new_n530), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n520), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n528), .B1(new_n527), .B2(new_n534), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT17), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT16), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(G1gat), .B1(new_n540), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(G8gat), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n541), .ZN(new_n548));
  INV_X1    g347(.A(G8gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n500), .A2(new_n502), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n520), .A2(new_n521), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT89), .B1(new_n555), .B2(new_n525), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n507), .A2(new_n518), .A3(new_n492), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n534), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n552), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n491), .B1(new_n537), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n553), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n551), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n553), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n565), .A3(new_n562), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n490), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g372(.A(KEYINPUT93), .B(new_n571), .C1(new_n560), .C2(new_n567), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n552), .B1(new_n535), .B2(new_n536), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n569), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n570), .B(KEYINPUT13), .Z(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n569), .A2(new_n570), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n560), .B2(new_n567), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(KEYINPUT18), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n489), .B1(new_n575), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n580), .ZN(new_n584));
  NOR3_X1   g383(.A1(new_n537), .A2(new_n559), .A3(new_n491), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n563), .B2(new_n566), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT18), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n587), .A2(new_n588), .B1(new_n577), .B2(new_n578), .ZN(new_n589));
  INV_X1    g388(.A(new_n489), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n589), .B(new_n590), .C1(new_n573), .C2(new_n574), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n583), .A2(KEYINPUT94), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n489), .C1(new_n575), .C2(new_n582), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n484), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G230gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n259), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT99), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT7), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT99), .B(new_n605), .C1(new_n599), .C2(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n599), .B2(new_n600), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G57gat), .B(G64gat), .Z(new_n614));
  AND2_X1   g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(KEYINPUT9), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G71gat), .B(G78gat), .Z(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n611), .A2(new_n619), .A3(new_n618), .A4(new_n612), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n598), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n623), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n598), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  OR2_X1    g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n627), .A2(new_n598), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n613), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n537), .A2(new_n561), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n564), .A2(new_n565), .A3(new_n638), .ZN(new_n640));
  NAND3_X1  g439(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  OR3_X1    g442(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n643), .B1(new_n639), .B2(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648));
  INV_X1    g447(.A(G232gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n259), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n647), .B(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n646), .A2(KEYINPUT100), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(KEYINPUT100), .Z(new_n653));
  AND2_X1   g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT21), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n552), .B1(new_n656), .B2(new_n620), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT95), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n658), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n620), .A2(new_n656), .ZN(new_n665));
  XNOR2_X1  g464(.A(G127gat), .B(G155gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT97), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(G183gat), .B(G211gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n664), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n596), .A2(new_n637), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n480), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n541), .ZN(G1324gat));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n429), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n549), .B2(new_n676), .ZN(new_n679));
  MUX2_X1   g478(.A(new_n678), .B(new_n679), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g479(.A(new_n476), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n286), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n673), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT101), .Z(G1326gat));
  INV_X1    g484(.A(new_n479), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n673), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n484), .ZN(new_n690));
  INV_X1    g489(.A(new_n671), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n636), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n595), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n655), .A3(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(G29gat), .A3(new_n480), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT45), .Z(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  INV_X1    g497(.A(new_n655), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n484), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n483), .A2(KEYINPUT102), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n472), .A2(new_n482), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n427), .A2(KEYINPUT103), .A3(new_n436), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT103), .B1(new_n427), .B2(new_n436), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n701), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n655), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n700), .B1(new_n707), .B2(new_n698), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n694), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n480), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(KEYINPUT104), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n710), .B2(KEYINPUT104), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n697), .B1(new_n711), .B2(new_n712), .ZN(G1328gat));
  NOR3_X1   g512(.A1(new_n695), .A2(G36gat), .A3(new_n429), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n709), .B2(new_n429), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  OAI21_X1  g516(.A(new_n494), .B1(new_n695), .B2(new_n286), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n476), .A2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n709), .B2(new_n458), .ZN(new_n722));
  OR3_X1    g521(.A1(new_n686), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT105), .B1(new_n686), .B2(G50gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n693), .A2(new_n699), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n596), .A2(new_n723), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n479), .A3(new_n694), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n730), .B2(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(KEYINPUT48), .B2(new_n731), .ZN(G1331gat));
  AND2_X1   g531(.A1(new_n672), .A2(new_n595), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n706), .A2(new_n636), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n480), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT106), .B(G57gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  INV_X1    g536(.A(new_n734), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT49), .B(G64gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n389), .A3(new_n739), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n734), .A2(new_n429), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT107), .Z(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n734), .B2(new_n681), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n286), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g546(.A1(new_n738), .A2(new_n479), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g548(.A1(new_n690), .A2(KEYINPUT44), .A3(new_n655), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n595), .A2(new_n671), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n636), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n437), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n427), .A2(KEYINPUT103), .A3(new_n436), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n472), .A2(new_n702), .A3(new_n482), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n702), .B1(new_n472), .B2(new_n482), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n699), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n750), .B(new_n755), .C1(new_n763), .C2(KEYINPUT44), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n480), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n704), .A2(new_n705), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n701), .A2(new_n703), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n655), .B(new_n753), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n655), .A4(new_n753), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n480), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n599), .A3(new_n636), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n765), .B1(new_n773), .B2(new_n775), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n389), .A2(new_n600), .A3(new_n636), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT109), .Z(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G92gat), .B1(new_n764), .B2(new_n429), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT44), .B1(new_n706), .B2(new_n655), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n783), .A2(new_n700), .A3(new_n754), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n600), .B1(new_n784), .B2(new_n389), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n768), .A2(KEYINPUT110), .A3(KEYINPUT51), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT51), .B1(new_n768), .B2(KEYINPUT110), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n789), .B2(new_n781), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n764), .B2(new_n681), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n424), .A2(new_n267), .A3(new_n636), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n773), .B2(new_n792), .ZN(G1338gat));
  NOR3_X1   g592(.A1(new_n458), .A2(G106gat), .A3(new_n637), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n786), .A2(new_n787), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n784), .B2(new_n479), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT53), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  OAI21_X1  g599(.A(G106gat), .B1(new_n764), .B2(new_n458), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT51), .B1(new_n763), .B2(new_n753), .ZN(new_n803));
  INV_X1    g602(.A(new_n771), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n794), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND4_X1   g604(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n772), .B2(new_n794), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n800), .B1(new_n807), .B2(new_n801), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(G1339gat));
  AND3_X1   g608(.A1(new_n672), .A2(new_n595), .A3(new_n637), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n577), .A2(new_n578), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n488), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n591), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n624), .A2(new_n625), .A3(new_n598), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n631), .B1(new_n626), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n635), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n820), .B2(new_n635), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n817), .B2(new_n819), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(new_n655), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n592), .A2(new_n594), .A3(new_n826), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n591), .A2(new_n636), .A3(new_n814), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n591), .A2(KEYINPUT113), .A3(new_n636), .A4(new_n814), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n828), .B1(new_n834), .B2(new_n699), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n811), .B1(new_n835), .B2(new_n691), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n480), .A2(new_n389), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n686), .A3(new_n424), .A4(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n595), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n592), .A2(new_n594), .A3(new_n826), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n832), .A2(new_n833), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n699), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n827), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n810), .B1(new_n847), .B2(new_n671), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n365), .A2(new_n425), .ZN(new_n849));
  NOR4_X1   g648(.A1(new_n848), .A2(new_n480), .A3(new_n389), .A4(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n595), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n244), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n843), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n242), .A3(new_n636), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n636), .A3(new_n841), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(G120gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n857), .B2(G120gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n842), .B2(new_n671), .ZN(new_n862));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n863), .A3(new_n691), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n842), .B2(new_n699), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n249), .A3(new_n655), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n681), .A2(new_n837), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n836), .B2(new_n364), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n821), .A2(new_n825), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n592), .A2(new_n594), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n655), .B1(new_n876), .B2(new_n830), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n671), .B1(new_n877), .B2(new_n828), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n874), .B(new_n686), .C1(new_n878), .C2(new_n811), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n872), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n595), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n681), .A2(new_n364), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n429), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n836), .A2(new_n774), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(G141gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n851), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n881), .B(new_n888), .C1(new_n891), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n896), .A3(new_n636), .ZN(new_n897));
  INV_X1    g696(.A(new_n880), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT59), .B(new_n896), .C1(new_n898), .C2(new_n636), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n686), .A2(KEYINPUT57), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n876), .A2(new_n830), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n699), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n827), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n877), .B2(new_n828), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n671), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(new_n811), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n874), .B1(new_n836), .B2(new_n364), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n636), .A3(new_n872), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n900), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n897), .B1(new_n899), .B2(new_n913), .ZN(G1345gat));
  NOR2_X1   g713(.A1(new_n671), .A2(new_n303), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n886), .A2(new_n691), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n898), .A2(new_n916), .B1(new_n303), .B2(new_n917), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n886), .B2(new_n655), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n699), .A2(new_n290), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n898), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n848), .A2(new_n774), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n849), .A2(new_n429), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n851), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n848), .A2(new_n479), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n774), .A2(new_n429), .A3(new_n286), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n223), .A3(new_n595), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n925), .A2(new_n929), .ZN(G1348gat));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n224), .A3(new_n637), .ZN(new_n931));
  AOI21_X1  g730(.A(G176gat), .B1(new_n924), .B2(new_n636), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n671), .A2(new_n211), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n922), .A2(new_n923), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n922), .A2(KEYINPUT122), .A3(new_n923), .A4(new_n936), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G183gat), .B1(new_n928), .B2(new_n671), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT60), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n945), .A2(KEYINPUT123), .A3(new_n946), .A4(new_n942), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n924), .A2(new_n231), .A3(new_n655), .ZN(new_n949));
  OAI21_X1  g748(.A(G190gat), .B1(new_n928), .B2(new_n699), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  NOR2_X1   g752(.A1(new_n882), .A2(new_n429), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n922), .A2(KEYINPUT124), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n836), .A2(new_n480), .A3(new_n954), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n851), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n774), .A2(new_n429), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n681), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n909), .A2(new_n910), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(G197gat), .A3(new_n851), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n960), .A2(new_n964), .ZN(G1352gat));
  INV_X1    g764(.A(new_n963), .ZN(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n966), .B2(new_n637), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n956), .A2(G204gat), .A3(new_n637), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1353gat));
  NAND2_X1  g769(.A1(new_n908), .A2(new_n811), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(new_n901), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT57), .B1(new_n848), .B2(new_n458), .ZN(new_n973));
  INV_X1    g772(.A(new_n962), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n972), .A2(new_n691), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g775(.A(G211gat), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT126), .B1(new_n963), .B2(new_n691), .ZN(new_n978));
  OAI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n963), .A2(KEYINPUT126), .A3(new_n691), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n975), .A2(new_n976), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(G211gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n671), .A2(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n955), .A2(new_n958), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n955), .A2(new_n987), .A3(new_n958), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n979), .A2(new_n983), .A3(new_n989), .ZN(G1354gat));
  NOR2_X1   g789(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n655), .B1(new_n963), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G218gat), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(G218gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n959), .A2(new_n995), .A3(new_n655), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1355gat));
endmodule


