

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753;

  INV_X1 U367 ( .A(n539), .ZN(n694) );
  OR2_X1 U368 ( .A1(n627), .A2(n606), .ZN(n440) );
  OR2_X1 U369 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X2 U370 ( .A1(n505), .A2(n500), .ZN(n648) );
  XNOR2_X2 U371 ( .A(G146), .B(n743), .ZN(n416) );
  OR2_X2 U372 ( .A1(n492), .A2(n692), .ZN(n539) );
  NOR2_X2 U373 ( .A1(G953), .A2(G237), .ZN(n471) );
  AND2_X1 U374 ( .A1(n506), .A2(n637), .ZN(n524) );
  OR2_X1 U375 ( .A1(n643), .A2(n516), .ZN(n522) );
  AND2_X1 U376 ( .A1(n648), .A2(n528), .ZN(n501) );
  AND2_X1 U377 ( .A1(n499), .A2(n596), .ZN(n505) );
  OR2_X1 U378 ( .A1(n498), .A2(n495), .ZN(n497) );
  XNOR2_X1 U379 ( .A(n515), .B(n514), .ZN(n726) );
  XNOR2_X1 U380 ( .A(n458), .B(KEYINPUT98), .ZN(n507) );
  AND2_X1 U381 ( .A1(n570), .A2(n569), .ZN(n597) );
  XNOR2_X1 U382 ( .A(n519), .B(KEYINPUT107), .ZN(n568) );
  XNOR2_X1 U383 ( .A(n440), .B(n439), .ZN(n545) );
  XNOR2_X1 U384 ( .A(n419), .B(n418), .ZN(n697) );
  XNOR2_X1 U385 ( .A(G146), .B(G125), .ZN(n429) );
  INV_X2 U386 ( .A(G953), .ZN(n427) );
  XNOR2_X1 U387 ( .A(G116), .B(G107), .ZN(n466) );
  XNOR2_X1 U388 ( .A(G119), .B(G113), .ZN(n410) );
  XNOR2_X1 U389 ( .A(G101), .B(KEYINPUT72), .ZN(n409) );
  XOR2_X1 U390 ( .A(KEYINPUT24), .B(KEYINPUT100), .Z(n390) );
  XNOR2_X1 U391 ( .A(G128), .B(KEYINPUT23), .ZN(n389) );
  NAND2_X1 U392 ( .A1(n364), .A2(KEYINPUT65), .ZN(n363) );
  INV_X1 U393 ( .A(n366), .ZN(n364) );
  XNOR2_X1 U394 ( .A(n470), .B(n469), .ZN(n517) );
  INV_X1 U395 ( .A(G478), .ZN(n469) );
  INV_X1 U396 ( .A(G902), .ZN(n481) );
  XNOR2_X1 U397 ( .A(n346), .B(n413), .ZN(n369) );
  AND2_X1 U398 ( .A1(n602), .A2(n601), .ZN(n746) );
  AND2_X1 U399 ( .A1(n524), .A2(n523), .ZN(n533) );
  AND2_X2 U400 ( .A1(n731), .A2(n746), .ZN(n674) );
  NAND2_X1 U401 ( .A1(n365), .A2(n361), .ZN(n360) );
  NAND2_X1 U402 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U403 ( .A1(n674), .A2(n352), .ZN(n365) );
  NAND2_X1 U404 ( .A1(n366), .A2(n353), .ZN(n362) );
  NOR2_X1 U405 ( .A1(n674), .A2(n359), .ZN(n358) );
  NAND2_X1 U406 ( .A1(n366), .A2(KEYINPUT65), .ZN(n359) );
  XNOR2_X1 U407 ( .A(G107), .B(G101), .ZN(n378) );
  XNOR2_X1 U408 ( .A(G116), .B(G137), .ZN(n414) );
  NOR2_X1 U409 ( .A1(n607), .A2(n351), .ZN(n366) );
  XNOR2_X1 U410 ( .A(G143), .B(G113), .ZN(n475) );
  XNOR2_X1 U411 ( .A(n482), .B(n345), .ZN(n518) );
  XNOR2_X1 U412 ( .A(G119), .B(G110), .ZN(n391) );
  XNOR2_X1 U413 ( .A(n462), .B(KEYINPUT106), .ZN(n463) );
  INV_X1 U414 ( .A(KEYINPUT22), .ZN(n489) );
  XNOR2_X1 U415 ( .A(n544), .B(n543), .ZN(n581) );
  AND2_X1 U416 ( .A1(n542), .A2(n541), .ZN(n544) );
  AND2_X1 U417 ( .A1(n652), .A2(n481), .ZN(n419) );
  OR2_X2 U418 ( .A1(n360), .A2(n358), .ZN(n611) );
  XNOR2_X1 U419 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U420 ( .A(n381), .B(n380), .ZN(n382) );
  INV_X1 U421 ( .A(KEYINPUT118), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n549), .B(KEYINPUT40), .ZN(n649) );
  XNOR2_X1 U423 ( .A(n572), .B(n370), .ZN(n573) );
  NAND2_X1 U424 ( .A1(n597), .A2(n571), .ZN(n572) );
  XNOR2_X1 U425 ( .A(n568), .B(n567), .ZN(n723) );
  XNOR2_X1 U426 ( .A(n354), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U427 ( .A1(n347), .A2(n355), .ZN(n354) );
  NAND2_X1 U428 ( .A1(n357), .A2(n356), .ZN(n355) );
  XOR2_X1 U429 ( .A(KEYINPUT13), .B(G475), .Z(n345) );
  XOR2_X1 U430 ( .A(n415), .B(n414), .Z(n346) );
  OR2_X1 U431 ( .A1(n716), .A2(n715), .ZN(n347) );
  XOR2_X1 U432 ( .A(n474), .B(KEYINPUT105), .Z(n348) );
  XOR2_X1 U433 ( .A(n464), .B(n463), .Z(n349) );
  XNOR2_X1 U434 ( .A(n548), .B(KEYINPUT39), .ZN(n594) );
  INV_X1 U435 ( .A(KEYINPUT65), .ZN(n367) );
  XOR2_X1 U436 ( .A(n561), .B(KEYINPUT64), .Z(n350) );
  AND2_X1 U437 ( .A1(n606), .A2(n603), .ZN(n351) );
  AND2_X1 U438 ( .A1(n606), .A2(n367), .ZN(n352) );
  OR2_X1 U439 ( .A1(n606), .A2(n367), .ZN(n353) );
  NAND2_X1 U440 ( .A1(n710), .A2(n709), .ZN(n357) );
  XNOR2_X1 U441 ( .A(n416), .B(n368), .ZN(n652) );
  XNOR2_X1 U442 ( .A(n369), .B(n426), .ZN(n368) );
  BUF_X1 U443 ( .A(n545), .Z(n599) );
  XNOR2_X2 U444 ( .A(n465), .B(n373), .ZN(n743) );
  XNOR2_X2 U445 ( .A(n431), .B(n372), .ZN(n465) );
  XOR2_X1 U446 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n370) );
  XOR2_X1 U447 ( .A(n390), .B(n389), .Z(n371) );
  INV_X1 U448 ( .A(KEYINPUT70), .ZN(n588) );
  XNOR2_X1 U449 ( .A(n562), .B(n350), .ZN(n591) );
  AND2_X1 U450 ( .A1(n492), .A2(n723), .ZN(n569) );
  INV_X1 U451 ( .A(KEYINPUT122), .ZN(n616) );
  XNOR2_X2 U452 ( .A(G143), .B(G128), .ZN(n431) );
  INV_X1 U453 ( .A(G134), .ZN(n372) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(G131), .ZN(n373) );
  INV_X1 U455 ( .A(G104), .ZN(n374) );
  NAND2_X1 U456 ( .A1(G110), .A2(n374), .ZN(n377) );
  INV_X1 U457 ( .A(G110), .ZN(n375) );
  NAND2_X1 U458 ( .A1(n375), .A2(G104), .ZN(n376) );
  NAND2_X1 U459 ( .A1(n377), .A2(n376), .ZN(n379) );
  XNOR2_X1 U460 ( .A(n379), .B(n378), .ZN(n383) );
  NAND2_X1 U461 ( .A1(G227), .A2(n427), .ZN(n381) );
  INV_X1 U462 ( .A(G140), .ZN(n380) );
  XOR2_X2 U463 ( .A(G137), .B(KEYINPUT68), .Z(n392) );
  INV_X1 U464 ( .A(KEYINPUT99), .ZN(n384) );
  XNOR2_X1 U465 ( .A(n392), .B(n384), .ZN(n744) );
  XNOR2_X1 U466 ( .A(n385), .B(n744), .ZN(n386) );
  XNOR2_X1 U467 ( .A(n416), .B(n386), .ZN(n664) );
  NAND2_X1 U468 ( .A1(n664), .A2(n481), .ZN(n388) );
  XOR2_X1 U469 ( .A(KEYINPUT71), .B(G469), .Z(n387) );
  XNOR2_X2 U470 ( .A(n388), .B(n387), .ZN(n553) );
  XNOR2_X2 U471 ( .A(n553), .B(KEYINPUT1), .ZN(n491) );
  XNOR2_X1 U472 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n371), .B(n393), .ZN(n396) );
  NAND2_X1 U474 ( .A1(G234), .A2(n427), .ZN(n394) );
  XOR2_X1 U475 ( .A(KEYINPUT8), .B(n394), .Z(n461) );
  NAND2_X1 U476 ( .A1(G221), .A2(n461), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n396), .B(n395), .ZN(n400) );
  XNOR2_X1 U478 ( .A(n429), .B(n380), .ZN(n398) );
  XOR2_X1 U479 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n397) );
  XNOR2_X1 U480 ( .A(n398), .B(n397), .ZN(n742) );
  INV_X1 U481 ( .A(n742), .ZN(n399) );
  XNOR2_X1 U482 ( .A(n400), .B(n399), .ZN(n659) );
  NAND2_X1 U483 ( .A1(n659), .A2(n481), .ZN(n405) );
  XNOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n401) );
  XNOR2_X1 U485 ( .A(n401), .B(G902), .ZN(n604) );
  NAND2_X1 U486 ( .A1(G234), .A2(n604), .ZN(n402) );
  XNOR2_X1 U487 ( .A(KEYINPUT20), .B(n402), .ZN(n406) );
  NAND2_X1 U488 ( .A1(G217), .A2(n406), .ZN(n403) );
  XNOR2_X1 U489 ( .A(n403), .B(KEYINPUT25), .ZN(n404) );
  XNOR2_X2 U490 ( .A(n405), .B(n404), .ZN(n492) );
  NAND2_X1 U491 ( .A1(G221), .A2(n406), .ZN(n407) );
  XNOR2_X1 U492 ( .A(n407), .B(KEYINPUT21), .ZN(n692) );
  NAND2_X1 U493 ( .A1(n491), .A2(n694), .ZN(n408) );
  XNOR2_X2 U494 ( .A(n408), .B(KEYINPUT76), .ZN(n512) );
  INV_X1 U495 ( .A(n512), .ZN(n420) );
  XNOR2_X1 U496 ( .A(n410), .B(n409), .ZN(n412) );
  XNOR2_X1 U497 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n411) );
  XNOR2_X1 U498 ( .A(n412), .B(n411), .ZN(n426) );
  NAND2_X1 U499 ( .A1(n471), .A2(G210), .ZN(n413) );
  XOR2_X1 U500 ( .A(KEYINPUT101), .B(KEYINPUT5), .Z(n415) );
  INV_X1 U501 ( .A(KEYINPUT102), .ZN(n417) );
  XOR2_X1 U502 ( .A(n417), .B(G472), .Z(n418) );
  XNOR2_X1 U503 ( .A(n697), .B(KEYINPUT6), .ZN(n566) );
  NAND2_X1 U504 ( .A1(n420), .A2(n566), .ZN(n421) );
  XNOR2_X2 U505 ( .A(n421), .B(KEYINPUT33), .ZN(n690) );
  XNOR2_X1 U506 ( .A(KEYINPUT16), .B(G110), .ZN(n422) );
  XNOR2_X1 U507 ( .A(n466), .B(n422), .ZN(n424) );
  INV_X1 U508 ( .A(G122), .ZN(n423) );
  XNOR2_X1 U509 ( .A(n423), .B(G104), .ZN(n477) );
  XNOR2_X1 U510 ( .A(n424), .B(n477), .ZN(n425) );
  XNOR2_X1 U511 ( .A(n426), .B(n425), .ZN(n737) );
  NAND2_X1 U512 ( .A1(n427), .A2(G224), .ZN(n428) );
  XNOR2_X1 U513 ( .A(n428), .B(KEYINPUT4), .ZN(n430) );
  XNOR2_X1 U514 ( .A(n430), .B(n429), .ZN(n434) );
  XNOR2_X1 U515 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n432) );
  XNOR2_X1 U516 ( .A(n431), .B(n432), .ZN(n433) );
  XNOR2_X1 U517 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U518 ( .A(n737), .B(n435), .ZN(n627) );
  INV_X1 U519 ( .A(n604), .ZN(n606) );
  INV_X1 U520 ( .A(G237), .ZN(n436) );
  NAND2_X1 U521 ( .A1(n436), .A2(n481), .ZN(n441) );
  NAND2_X1 U522 ( .A1(n441), .A2(G210), .ZN(n438) );
  INV_X1 U523 ( .A(KEYINPUT79), .ZN(n437) );
  XNOR2_X1 U524 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U525 ( .A1(n441), .A2(G214), .ZN(n442) );
  XNOR2_X1 U526 ( .A(n442), .B(KEYINPUT94), .ZN(n564) );
  INV_X1 U527 ( .A(n564), .ZN(n683) );
  OR2_X2 U528 ( .A1(n545), .A2(n683), .ZN(n443) );
  XNOR2_X2 U529 ( .A(n443), .B(KEYINPUT19), .ZN(n574) );
  XOR2_X1 U530 ( .A(KEYINPUT95), .B(KEYINPUT14), .Z(n445) );
  NAND2_X1 U531 ( .A1(G237), .A2(G234), .ZN(n444) );
  XNOR2_X1 U532 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U533 ( .A(KEYINPUT74), .B(n446), .ZN(n450) );
  NAND2_X1 U534 ( .A1(n450), .A2(G952), .ZN(n448) );
  INV_X1 U535 ( .A(KEYINPUT96), .ZN(n447) );
  XNOR2_X1 U536 ( .A(n448), .B(n447), .ZN(n711) );
  AND2_X1 U537 ( .A1(n711), .A2(n427), .ZN(n708) );
  AND2_X1 U538 ( .A1(G953), .A2(G902), .ZN(n449) );
  NAND2_X1 U539 ( .A1(n450), .A2(n449), .ZN(n536) );
  NOR2_X1 U540 ( .A1(G898), .A2(n536), .ZN(n451) );
  NOR2_X1 U541 ( .A1(n708), .A2(n451), .ZN(n452) );
  XNOR2_X1 U542 ( .A(n452), .B(KEYINPUT97), .ZN(n453) );
  NAND2_X1 U543 ( .A1(n574), .A2(n453), .ZN(n457) );
  XNOR2_X1 U544 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n455) );
  INV_X1 U545 ( .A(KEYINPUT66), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U547 ( .A(n457), .B(n456), .ZN(n513) );
  INV_X1 U548 ( .A(n513), .ZN(n458) );
  NAND2_X1 U549 ( .A1(n690), .A2(n507), .ZN(n460) );
  XNOR2_X1 U550 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n459) );
  XNOR2_X1 U551 ( .A(n460), .B(n459), .ZN(n484) );
  NAND2_X1 U552 ( .A1(G217), .A2(n461), .ZN(n464) );
  XOR2_X1 U553 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n462) );
  XNOR2_X1 U554 ( .A(n466), .B(G122), .ZN(n467) );
  XNOR2_X1 U555 ( .A(n465), .B(n467), .ZN(n468) );
  XNOR2_X1 U556 ( .A(n349), .B(n468), .ZN(n612) );
  NAND2_X1 U557 ( .A1(n612), .A2(n481), .ZN(n470) );
  INV_X1 U558 ( .A(n517), .ZN(n521) );
  XOR2_X1 U559 ( .A(KEYINPUT12), .B(KEYINPUT104), .Z(n473) );
  NAND2_X1 U560 ( .A1(n471), .A2(G214), .ZN(n472) );
  XNOR2_X1 U561 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U562 ( .A(G131), .B(KEYINPUT11), .Z(n476) );
  XNOR2_X1 U563 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U564 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U565 ( .A(n348), .B(n479), .ZN(n480) );
  XNOR2_X1 U566 ( .A(n480), .B(n742), .ZN(n618) );
  NAND2_X1 U567 ( .A1(n618), .A2(n481), .ZN(n482) );
  NAND2_X1 U568 ( .A1(n521), .A2(n518), .ZN(n579) );
  INV_X1 U569 ( .A(n579), .ZN(n483) );
  NAND2_X1 U570 ( .A1(n484), .A2(n483), .ZN(n486) );
  INV_X1 U571 ( .A(KEYINPUT35), .ZN(n485) );
  XNOR2_X2 U572 ( .A(n486), .B(n485), .ZN(n650) );
  INV_X1 U573 ( .A(n518), .ZN(n520) );
  AND2_X1 U574 ( .A1(n520), .A2(n517), .ZN(n681) );
  INV_X1 U575 ( .A(n692), .ZN(n487) );
  NAND2_X1 U576 ( .A1(n681), .A2(n487), .ZN(n488) );
  NOR2_X1 U577 ( .A1(n513), .A2(n488), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n490), .B(n489), .ZN(n498) );
  NAND2_X1 U579 ( .A1(n491), .A2(n492), .ZN(n493) );
  XNOR2_X1 U580 ( .A(n493), .B(KEYINPUT108), .ZN(n494) );
  OR2_X1 U581 ( .A1(n494), .A2(n566), .ZN(n495) );
  XNOR2_X1 U582 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n496) );
  XNOR2_X2 U583 ( .A(n497), .B(n496), .ZN(n647) );
  INV_X1 U584 ( .A(n498), .ZN(n499) );
  INV_X1 U585 ( .A(n491), .ZN(n596) );
  AND2_X1 U586 ( .A1(n697), .A2(n492), .ZN(n500) );
  INV_X1 U587 ( .A(KEYINPUT44), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n647), .A2(n501), .ZN(n502) );
  INV_X1 U589 ( .A(KEYINPUT85), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n502), .A2(n529), .ZN(n503) );
  NAND2_X1 U591 ( .A1(n650), .A2(n503), .ZN(n506) );
  NOR2_X1 U592 ( .A1(n566), .A2(n492), .ZN(n504) );
  NAND2_X1 U593 ( .A1(n505), .A2(n504), .ZN(n637) );
  INV_X1 U594 ( .A(n507), .ZN(n510) );
  AND2_X1 U595 ( .A1(n697), .A2(n694), .ZN(n508) );
  NAND2_X1 U596 ( .A1(n508), .A2(n553), .ZN(n509) );
  OR2_X1 U597 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U598 ( .A(n511), .B(KEYINPUT103), .ZN(n643) );
  OR2_X1 U599 ( .A1(n697), .A2(n512), .ZN(n691) );
  OR2_X1 U600 ( .A1(n513), .A2(n691), .ZN(n515) );
  INV_X1 U601 ( .A(KEYINPUT31), .ZN(n514) );
  INV_X1 U602 ( .A(n726), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U604 ( .A1(n521), .A2(n520), .ZN(n727) );
  INV_X1 U605 ( .A(n727), .ZN(n717) );
  OR2_X1 U606 ( .A1(n568), .A2(n717), .ZN(n686) );
  XNOR2_X1 U607 ( .A(n686), .B(KEYINPUT82), .ZN(n576) );
  NAND2_X1 U608 ( .A1(n522), .A2(n576), .ZN(n523) );
  OR2_X1 U609 ( .A1(n650), .A2(KEYINPUT85), .ZN(n527) );
  AND2_X1 U610 ( .A1(n648), .A2(KEYINPUT44), .ZN(n525) );
  AND2_X1 U611 ( .A1(n525), .A2(n647), .ZN(n526) );
  NAND2_X1 U612 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U613 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U614 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U615 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U616 ( .A(n534), .B(KEYINPUT45), .ZN(n731) );
  NOR2_X1 U617 ( .A1(n697), .A2(n683), .ZN(n535) );
  XNOR2_X1 U618 ( .A(n535), .B(KEYINPUT30), .ZN(n542) );
  XNOR2_X1 U619 ( .A(KEYINPUT110), .B(n536), .ZN(n537) );
  NOR2_X1 U620 ( .A1(G900), .A2(n537), .ZN(n538) );
  NOR2_X1 U621 ( .A1(n708), .A2(n538), .ZN(n550) );
  NOR2_X1 U622 ( .A1(n539), .A2(n550), .ZN(n540) );
  AND2_X1 U623 ( .A1(n553), .A2(n540), .ZN(n541) );
  INV_X1 U624 ( .A(KEYINPUT77), .ZN(n543) );
  INV_X1 U625 ( .A(KEYINPUT75), .ZN(n546) );
  XNOR2_X1 U626 ( .A(n546), .B(KEYINPUT38), .ZN(n547) );
  XNOR2_X1 U627 ( .A(n599), .B(n547), .ZN(n555) );
  NAND2_X1 U628 ( .A1(n581), .A2(n555), .ZN(n548) );
  NAND2_X1 U629 ( .A1(n594), .A2(n568), .ZN(n549) );
  NOR2_X1 U630 ( .A1(n692), .A2(n550), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n492), .A2(n563), .ZN(n551) );
  NOR2_X1 U632 ( .A1(n697), .A2(n551), .ZN(n552) );
  XNOR2_X1 U633 ( .A(n552), .B(KEYINPUT28), .ZN(n554) );
  AND2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n681), .A2(n564), .ZN(n556) );
  INV_X1 U636 ( .A(n555), .ZN(n684) );
  OR2_X1 U637 ( .A1(n556), .A2(n684), .ZN(n559) );
  INV_X1 U638 ( .A(KEYINPUT111), .ZN(n557) );
  XNOR2_X1 U639 ( .A(n557), .B(KEYINPUT41), .ZN(n558) );
  XNOR2_X1 U640 ( .A(n559), .B(n558), .ZN(n703) );
  NAND2_X1 U641 ( .A1(n575), .A2(n703), .ZN(n560) );
  XNOR2_X1 U642 ( .A(n560), .B(KEYINPUT42), .ZN(n635) );
  NAND2_X1 U643 ( .A1(n649), .A2(n635), .ZN(n562) );
  XNOR2_X1 U644 ( .A(KEYINPUT84), .B(KEYINPUT46), .ZN(n561) );
  AND2_X1 U645 ( .A1(n564), .A2(n563), .ZN(n565) );
  AND2_X1 U646 ( .A1(n566), .A2(n565), .ZN(n570) );
  INV_X1 U647 ( .A(KEYINPUT109), .ZN(n567) );
  INV_X1 U648 ( .A(n599), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n573), .A2(n491), .ZN(n730) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n582), .A2(KEYINPUT47), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n578) );
  AND2_X1 U653 ( .A1(n730), .A2(n578), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n579), .A2(n599), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n722) );
  INV_X1 U656 ( .A(n582), .ZN(n718) );
  NAND2_X1 U657 ( .A1(n718), .A2(n686), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n583), .A2(KEYINPUT47), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n722), .A2(n584), .ZN(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT81), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U664 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n593), .B(n592), .ZN(n602) );
  INV_X1 U666 ( .A(n594), .ZN(n595) );
  OR2_X1 U667 ( .A1(n595), .A2(n727), .ZN(n640) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT43), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n638) );
  AND2_X1 U671 ( .A1(n640), .A2(n638), .ZN(n601) );
  INV_X1 U672 ( .A(KEYINPUT2), .ZN(n608) );
  NOR2_X1 U673 ( .A1(n608), .A2(KEYINPUT83), .ZN(n603) );
  NAND2_X1 U674 ( .A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n607) );
  INV_X1 U676 ( .A(n674), .ZN(n609) );
  OR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n610) );
  AND2_X2 U678 ( .A1(n611), .A2(n610), .ZN(n663) );
  NAND2_X1 U679 ( .A1(n663), .A2(G478), .ZN(n613) );
  XNOR2_X1 U680 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U681 ( .A(G952), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n614), .A2(G953), .ZN(n670) );
  NAND2_X1 U683 ( .A1(n615), .A2(n670), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n617), .B(n616), .ZN(G63) );
  NAND2_X1 U685 ( .A1(n663), .A2(G475), .ZN(n620) );
  XOR2_X1 U686 ( .A(n618), .B(KEYINPUT59), .Z(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U688 ( .A1(n621), .A2(n670), .ZN(n623) );
  INV_X1 U689 ( .A(KEYINPUT60), .ZN(n622) );
  XNOR2_X1 U690 ( .A(n623), .B(n622), .ZN(G60) );
  NAND2_X1 U691 ( .A1(n663), .A2(G210), .ZN(n629) );
  XOR2_X1 U692 ( .A(KEYINPUT88), .B(KEYINPUT54), .Z(n625) );
  XNOR2_X1 U693 ( .A(KEYINPUT55), .B(KEYINPUT87), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U697 ( .A1(n630), .A2(n670), .ZN(n632) );
  INV_X1 U698 ( .A(KEYINPUT56), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(G51) );
  NAND2_X1 U700 ( .A1(n718), .A2(n723), .ZN(n634) );
  XOR2_X1 U701 ( .A(G146), .B(KEYINPUT115), .Z(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G48) );
  XNOR2_X1 U703 ( .A(G137), .B(KEYINPUT127), .ZN(n636) );
  XOR2_X1 U704 ( .A(n636), .B(n635), .Z(G39) );
  XNOR2_X1 U705 ( .A(n637), .B(G101), .ZN(G3) );
  XNOR2_X1 U706 ( .A(n638), .B(G140), .ZN(G42) );
  NAND2_X1 U707 ( .A1(n643), .A2(n723), .ZN(n639) );
  XNOR2_X1 U708 ( .A(n639), .B(G104), .ZN(G6) );
  XNOR2_X1 U709 ( .A(n640), .B(G134), .ZN(G36) );
  XOR2_X1 U710 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n642) );
  XNOR2_X1 U711 ( .A(G107), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n643), .A2(n717), .ZN(n644) );
  XOR2_X1 U714 ( .A(n645), .B(n644), .Z(G9) );
  XNOR2_X1 U715 ( .A(G119), .B(KEYINPUT126), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G21) );
  XNOR2_X1 U717 ( .A(n648), .B(G110), .ZN(G12) );
  XNOR2_X1 U718 ( .A(n649), .B(G131), .ZN(G33) );
  XNOR2_X1 U719 ( .A(n650), .B(G122), .ZN(G24) );
  NAND2_X1 U720 ( .A1(n663), .A2(G472), .ZN(n654) );
  XNOR2_X1 U721 ( .A(KEYINPUT90), .B(KEYINPUT62), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(n670), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT86), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n658), .B(n657), .ZN(G57) );
  NAND2_X1 U728 ( .A1(n663), .A2(G217), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n661), .A2(n670), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U732 ( .A1(n663), .A2(G469), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n666) );
  XNOR2_X1 U734 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n664), .B(n667), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n669), .B(n668), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT121), .ZN(G54) );
  INV_X1 U740 ( .A(KEYINPUT80), .ZN(n673) );
  XNOR2_X1 U741 ( .A(n675), .B(KEYINPUT2), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n690), .A2(n703), .ZN(n677) );
  INV_X1 U743 ( .A(KEYINPUT117), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n716) );
  NAND2_X1 U746 ( .A1(n716), .A2(n427), .ZN(n710) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT116), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n706) );
  INV_X1 U754 ( .A(n691), .ZN(n701) );
  NAND2_X1 U755 ( .A1(n692), .A2(n492), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n693), .B(KEYINPUT49), .ZN(n699) );
  NOR2_X1 U757 ( .A1(n694), .A2(n491), .ZN(n695) );
  XOR2_X1 U758 ( .A(KEYINPUT50), .B(n695), .Z(n696) );
  NAND2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U762 ( .A(n702), .B(KEYINPUT51), .ZN(n704) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U765 ( .A(n707), .B(KEYINPUT52), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n712), .A2(n708), .ZN(n709) );
  NAND2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n714) );
  AND2_X1 U768 ( .A1(n427), .A2(KEYINPUT118), .ZN(n713) );
  NAND2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n720) );
  XOR2_X1 U771 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n719) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U773 ( .A(G128), .B(n721), .ZN(G30) );
  XNOR2_X1 U774 ( .A(G143), .B(n722), .ZN(G45) );
  INV_X1 U775 ( .A(n723), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n724), .A2(n726), .ZN(n725) );
  XOR2_X1 U777 ( .A(G113), .B(n725), .Z(G15) );
  NOR2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U779 ( .A(G116), .B(n728), .Z(G18) );
  XOR2_X1 U780 ( .A(G125), .B(KEYINPUT37), .Z(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(n729), .ZN(G27) );
  AND2_X1 U782 ( .A1(n731), .A2(n427), .ZN(n736) );
  INV_X1 U783 ( .A(G898), .ZN(n734) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n732) );
  XOR2_X1 U785 ( .A(KEYINPUT61), .B(n732), .Z(n733) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n741) );
  XNOR2_X1 U788 ( .A(n737), .B(KEYINPUT124), .ZN(n739) );
  NOR2_X1 U789 ( .A1(n427), .A2(G898), .ZN(n738) );
  NOR2_X1 U790 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U791 ( .A(n741), .B(n740), .Z(G69) );
  XOR2_X1 U792 ( .A(n743), .B(n742), .Z(n745) );
  XOR2_X1 U793 ( .A(n745), .B(n744), .Z(n748) );
  XOR2_X1 U794 ( .A(n746), .B(n748), .Z(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(n427), .ZN(n753) );
  XNOR2_X1 U796 ( .A(G227), .B(n748), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(G900), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT125), .B(n750), .Z(n751) );
  NAND2_X1 U799 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(G72) );
endmodule

