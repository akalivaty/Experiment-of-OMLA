//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n451, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g025(.A(G2106), .ZN(new_n451));
  NOR2_X1   g026(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XNOR2_X1  g034(.A(new_n458), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n455), .A2(new_n451), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT68), .Z(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G137), .A4(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  INV_X1    g048(.A(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n464), .B1(new_n474), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n470), .A2(new_n498), .A3(G138), .A4(new_n464), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT70), .B(G88), .Z(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n505), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT71), .Z(new_n518));
  AOI21_X1  g093(.A(new_n506), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n505), .A2(new_n510), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n522), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n502), .A2(new_n504), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n534), .B1(new_n535), .B2(new_n513), .C1(new_n536), .C2(new_n511), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n511), .A2(new_n539), .B1(new_n513), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n506), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  NAND4_X1  g125(.A1(new_n507), .A2(new_n509), .A3(G53), .A4(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n505), .A2(new_n510), .A3(G91), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n531), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(G299));
  INV_X1    g133(.A(G166), .ZN(G303));
  OAI21_X1  g134(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n561));
  INV_X1    g136(.A(G87), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n511), .ZN(G288));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n511), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n502), .A2(new_n504), .A3(G61), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT72), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n506), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n564), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n523), .A2(G86), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n570), .B(KEYINPUT72), .Z(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n575), .B2(new_n568), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT73), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G305));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  INV_X1    g154(.A(G47), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n511), .A2(new_n579), .B1(new_n513), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n506), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n511), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n531), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n587), .A2(new_n590), .B1(G651), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n521), .A2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n586), .B1(new_n597), .B2(G868), .ZN(G321));
  XOR2_X1   g173(.A(G321), .B(KEYINPUT74), .Z(G284));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NOR2_X1   g180(.A1(new_n596), .A2(G559), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n544), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(KEYINPUT75), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(KEYINPUT75), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n484), .A2(G135), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n484), .A2(KEYINPUT77), .A3(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n482), .A2(G123), .ZN(new_n619));
  AND4_X1   g194(.A1(new_n614), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n484), .A2(G2104), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT13), .B(G2100), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT79), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT78), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n639), .B(new_n640), .Z(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(G14), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n645), .B2(new_n646), .ZN(new_n652));
  AOI21_X1  g227(.A(KEYINPUT18), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(KEYINPUT20), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(KEYINPUT20), .C2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G27), .ZN(new_n675));
  OAI21_X1  g250(.A(KEYINPUT94), .B1(new_n675), .B2(G29), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n675), .A2(KEYINPUT94), .A3(G29), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n677), .C1(G164), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2078), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n484), .A2(G139), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT25), .Z(new_n683));
  AOI22_X1  g258(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT90), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n681), .B(new_n683), .C1(new_n685), .C2(new_n464), .ZN(new_n686));
  MUX2_X1   g261(.A(G33), .B(new_n686), .S(G29), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  INV_X1    g263(.A(G2072), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n678), .A2(G26), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n482), .A2(G128), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n484), .A2(G140), .ZN(new_n694));
  NOR2_X1   g269(.A1(G104), .A2(G2105), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n692), .B1(new_n697), .B2(G29), .ZN(new_n698));
  MUX2_X1   g273(.A(new_n692), .B(new_n698), .S(KEYINPUT28), .Z(new_n699));
  INV_X1    g274(.A(G2067), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(KEYINPUT24), .A2(G34), .ZN(new_n702));
  NOR2_X1   g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n702), .A2(new_n703), .A3(G29), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n480), .B2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G2084), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR4_X1   g282(.A1(new_n690), .A2(new_n691), .A3(new_n701), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT93), .B1(G5), .B2(G16), .ZN(new_n709));
  OR3_X1    g284(.A1(KEYINPUT93), .A2(G5), .A3(G16), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n710), .C1(G301), .C2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n620), .A2(G29), .ZN(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n716), .A2(KEYINPUT92), .A3(KEYINPUT30), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT92), .B1(new_n716), .B2(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n678), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n717), .B(new_n719), .C1(KEYINPUT30), .C2(new_n716), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n714), .A2(new_n715), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  OR2_X1    g297(.A1(G29), .A2(G32), .ZN(new_n723));
  AOI22_X1  g298(.A1(G129), .A2(new_n482), .B1(new_n484), .B2(G141), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n678), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n712), .A2(new_n713), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n711), .A2(G4), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n596), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1348), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n711), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n711), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n734), .A2(new_n735), .B1(new_n737), .B2(G1966), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n721), .A2(new_n722), .A3(new_n731), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n678), .A2(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n678), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G2090), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n729), .B2(new_n730), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n544), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n737), .A2(G1966), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n739), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G299), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT23), .B1(new_n750), .B2(new_n711), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n711), .A2(G20), .ZN(new_n752));
  MUX2_X1   g327(.A(KEYINPUT23), .B(new_n751), .S(new_n752), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT96), .B(G1956), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n753), .B(new_n754), .Z(new_n755));
  NOR2_X1   g330(.A1(new_n742), .A2(G2090), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(KEYINPUT95), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(KEYINPUT95), .ZN(new_n758));
  INV_X1    g333(.A(new_n734), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(G1348), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n708), .A2(new_n749), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n484), .A2(G131), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT83), .ZN(new_n764));
  OR2_X1    g339(.A1(G95), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n482), .A2(G119), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT84), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n764), .A2(new_n770), .A3(new_n766), .A4(new_n767), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n678), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n678), .A2(G25), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT35), .B(G1991), .ZN(new_n775));
  OR3_X1    g350(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n772), .B2(new_n774), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n711), .A2(G23), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G288), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(KEYINPUT33), .B(new_n779), .C1(G288), .C2(G16), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1976), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n780), .A2(new_n781), .ZN(new_n787));
  OAI21_X1  g362(.A(G1976), .B1(new_n787), .B2(new_n783), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n711), .A2(G6), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G305), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT32), .B(G1981), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT87), .Z(new_n793));
  OR2_X1    g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(G16), .B1(new_n515), .B2(new_n519), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n711), .A2(G22), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n791), .B2(new_n793), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n789), .A2(new_n794), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n778), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G24), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT85), .B1(new_n805), .B2(G16), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n805), .A2(KEYINPUT85), .A3(G16), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n806), .B(new_n807), .C1(new_n584), .C2(new_n711), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT86), .B(G1986), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(KEYINPUT88), .B1(new_n801), .B2(KEYINPUT34), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n801), .A2(KEYINPUT88), .A3(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n804), .B(new_n810), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(KEYINPUT89), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n777), .B(new_n776), .C1(new_n801), .C2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n820), .B2(new_n812), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n816), .B1(new_n821), .B2(new_n810), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n762), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n814), .A2(KEYINPUT89), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n816), .A3(new_n810), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT36), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n680), .B(new_n761), .C1(new_n823), .C2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n826), .ZN(new_n828));
  INV_X1    g403(.A(new_n680), .ZN(new_n829));
  INV_X1    g404(.A(new_n761), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G150));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT98), .B(G55), .Z(new_n833));
  OAI22_X1  g408(.A1(new_n511), .A2(new_n832), .B1(new_n513), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n505), .A2(G67), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n506), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G860), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n834), .A2(new_n837), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n544), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT99), .B1(new_n834), .B2(new_n837), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n544), .A2(new_n840), .A3(new_n841), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n596), .A2(new_n604), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n839), .B1(new_n852), .B2(G860), .ZN(G145));
  XNOR2_X1  g428(.A(new_n488), .B(KEYINPUT100), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n620), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n769), .A2(new_n771), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n482), .A2(G130), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n484), .A2(G142), .ZN(new_n862));
  NOR2_X1   g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n624), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n865), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n860), .A3(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n859), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n858), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n728), .B(new_n697), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(new_n686), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n686), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n497), .A2(new_n499), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n490), .A2(KEYINPUT101), .A3(new_n494), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT101), .B1(new_n490), .B2(new_n494), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n495), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n879), .A2(new_n886), .A3(new_n880), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n876), .B2(new_n877), .ZN(new_n888));
  AND4_X1   g463(.A1(KEYINPUT104), .A2(new_n874), .A3(new_n884), .A4(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(KEYINPUT104), .A2(new_n874), .B1(new_n884), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n857), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT105), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(new_n857), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  AND4_X1   g471(.A1(new_n884), .A2(new_n888), .A3(new_n871), .A4(new_n873), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n884), .A2(new_n888), .B1(new_n871), .B2(new_n873), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n856), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT103), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(new_n856), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT40), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n895), .A2(new_n903), .A3(new_n906), .A4(new_n896), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(G395));
  XOR2_X1   g483(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n847), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n606), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n847), .B(KEYINPUT106), .ZN(new_n913));
  INV_X1    g488(.A(new_n606), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n597), .A2(new_n750), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n596), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n921), .A3(new_n917), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n596), .A2(G299), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n750), .B1(new_n595), .B2(new_n594), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT41), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n912), .B2(new_n915), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n909), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n909), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n912), .A2(new_n915), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n929), .B(new_n919), .C1(new_n930), .C2(new_n926), .ZN(new_n931));
  INV_X1    g506(.A(G288), .ZN(new_n932));
  NAND2_X1  g507(.A1(G290), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n584), .A2(G288), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G303), .B1(new_n573), .B2(new_n577), .ZN(new_n936));
  NOR2_X1   g511(.A1(G305), .A2(G166), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT107), .B1(new_n933), .B2(new_n934), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n936), .A2(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n928), .A2(new_n931), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n928), .B2(new_n931), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G868), .B2(new_n840), .ZN(G295));
  OAI21_X1  g523(.A(new_n947), .B1(G868), .B2(new_n840), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  INV_X1    g526(.A(new_n918), .ZN(new_n952));
  XNOR2_X1  g527(.A(G286), .B(G301), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n846), .B2(new_n845), .ZN(new_n954));
  NAND2_X1  g529(.A1(G168), .A2(G301), .ZN(new_n955));
  NAND2_X1  g530(.A1(G171), .A2(G286), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n847), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n918), .A2(new_n963), .A3(KEYINPUT41), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n953), .A2(new_n846), .A3(new_n845), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n847), .A2(new_n957), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n952), .B(KEYINPUT110), .C1(new_n954), .C2(new_n958), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n961), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n944), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n926), .A2(new_n965), .A3(new_n966), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n943), .A3(new_n959), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(new_n896), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n951), .B1(new_n974), .B2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n896), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n943), .B1(new_n971), .B2(new_n959), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(KEYINPUT43), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n950), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n970), .B2(new_n973), .ZN(new_n982));
  NOR4_X1   g557(.A1(new_n982), .A2(new_n978), .A3(KEYINPUT111), .A4(new_n951), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n970), .A2(new_n973), .A3(new_n981), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI22_X1  g561(.A1(new_n980), .A2(new_n983), .B1(KEYINPUT44), .B2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n887), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n472), .A2(new_n478), .A3(G40), .A4(new_n479), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n995));
  NAND2_X1  g570(.A1(G290), .A2(G1986), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n995), .B(new_n996), .Z(new_n997));
  NOR2_X1   g572(.A1(new_n858), .A2(new_n775), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n858), .A2(new_n775), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n728), .B(G1996), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n697), .B(G2067), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n993), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n887), .A2(new_n1006), .A3(new_n988), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n991), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  INV_X1    g586(.A(new_n495), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n879), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n988), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n990), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n1008), .A4(new_n1007), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G164), .B2(G1384), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n991), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n796), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1011), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G166), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1027), .A2(KEYINPUT55), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1011), .A2(new_n1017), .A3(new_n1022), .A4(KEYINPUT114), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1025), .A2(G8), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1033), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1022), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n991), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1006), .B1(new_n887), .B2(new_n988), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(G2090), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n574), .A2(new_n565), .A3(new_n576), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1043), .A2(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(G1981), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n887), .A2(new_n988), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n990), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n1026), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n785), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(G8), .C1(new_n1049), .C2(new_n990), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT52), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1058), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n785), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1051), .A2(new_n1060), .A3(new_n1056), .A4(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1053), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1035), .A2(new_n1042), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1007), .A2(new_n706), .A3(new_n991), .A4(new_n1009), .ZN(new_n1065));
  NOR3_X1   g640(.A1(G164), .A2(new_n1019), .A3(G1384), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n989), .A2(new_n1066), .A3(new_n990), .ZN(new_n1067));
  OAI211_X1 g642(.A(G168), .B(new_n1065), .C1(new_n1067), .C2(G1966), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(G8), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT122), .A3(KEYINPUT51), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1067), .B2(G1966), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1072), .A2(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G286), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1068), .A2(new_n1078), .A3(G8), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1064), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(G1996), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1018), .A2(new_n1082), .A3(new_n991), .A4(new_n1020), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n990), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT119), .A3(new_n1082), .A4(new_n1018), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1049), .B2(new_n990), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n544), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1093), .A3(new_n544), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1007), .A2(new_n991), .A3(new_n1009), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1096), .A2(new_n735), .B1(new_n1050), .B2(new_n700), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1097), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n596), .B1(new_n1097), .B2(KEYINPUT60), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1098), .A2(new_n1099), .B1(KEYINPUT60), .B2(new_n1097), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(G299), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(G299), .A2(new_n1101), .A3(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1049), .A2(KEYINPUT50), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1384), .B1(new_n879), .B2(new_n1012), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n990), .B1(new_n1006), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1956), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n1018), .A2(new_n991), .A3(new_n1020), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1105), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1956), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1114));
  AND3_X1   g689(.A1(G299), .A2(new_n1101), .A3(KEYINPUT57), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1102), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1086), .A2(new_n1018), .A3(new_n1110), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1112), .A2(new_n1118), .A3(new_n1119), .A4(KEYINPUT61), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(KEYINPUT61), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(KEYINPUT61), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1095), .A2(new_n1100), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1112), .B1(new_n596), .B2(new_n1097), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1384), .B1(new_n883), .B2(new_n879), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT124), .B(new_n991), .C1(new_n1130), .C2(KEYINPUT45), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n989), .B2(new_n990), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(G2078), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(new_n1018), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G2078), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1018), .A2(new_n1137), .A3(new_n991), .A4(new_n1020), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT123), .B(G1961), .Z(new_n1139));
  AOI22_X1  g714(.A1(new_n1134), .A2(new_n1138), .B1(new_n1096), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1129), .B1(new_n1142), .B2(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1067), .A2(new_n1135), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(G301), .A3(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1145), .C1(KEYINPUT126), .C2(new_n1142), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1136), .A2(new_n1140), .A3(G301), .ZN(new_n1147));
  AOI21_X1  g722(.A(G301), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1129), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT125), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n1129), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1081), .A2(new_n1128), .A3(new_n1146), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1025), .A2(G8), .A3(new_n1034), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1036), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1072), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1035), .A3(new_n1063), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1073), .A2(G168), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1064), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1157), .B1(new_n1155), .B2(new_n1036), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1165), .A2(KEYINPUT117), .A3(new_n1035), .A4(new_n1063), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1035), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1053), .A2(new_n785), .A3(new_n932), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1044), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1168), .A2(new_n1063), .B1(new_n1170), .B2(new_n1051), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1154), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1079), .A2(new_n1077), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1074), .B(new_n1071), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1175), .A2(new_n1176), .A3(KEYINPUT62), .ZN(new_n1177));
  AND4_X1   g752(.A1(new_n1035), .A2(new_n1063), .A3(new_n1148), .A4(new_n1042), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1175), .B2(KEYINPUT62), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1176), .B1(new_n1175), .B2(KEYINPUT62), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1005), .B1(new_n1172), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n998), .A2(new_n1003), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n697), .A2(G2067), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n992), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n993), .B1(new_n728), .B2(new_n1002), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n993), .A2(KEYINPUT46), .A3(new_n1082), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT46), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n992), .B2(G1996), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT47), .Z(new_n1191));
  NAND2_X1  g766(.A1(new_n1004), .A2(new_n993), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n993), .A2(new_n994), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1185), .B(new_n1191), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1182), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(G319), .ZN(new_n1198));
  AOI211_X1 g772(.A(new_n1198), .B(G227), .C1(new_n984), .C2(new_n985), .ZN(new_n1199));
  NOR2_X1   g773(.A1(G401), .A2(G229), .ZN(new_n1200));
  AND3_X1   g774(.A1(new_n1199), .A2(new_n904), .A3(new_n1200), .ZN(G308));
  NAND3_X1  g775(.A1(new_n1199), .A2(new_n904), .A3(new_n1200), .ZN(G225));
endmodule


