//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  NAND2_X1  g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n203), .A2(KEYINPUT22), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(KEYINPUT73), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n203), .A2(new_n204), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n206), .A2(new_n207), .B1(new_n212), .B2(new_n202), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G226gat), .ZN(new_n217));
  INV_X1    g016(.A(G233gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n223), .B(new_n224), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT27), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n228), .A3(new_n224), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n229), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT66), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n226), .A2(new_n230), .A3(new_n233), .A4(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  INV_X1    g048(.A(G169gat), .ZN(new_n250));
  INV_X1    g049(.A(G176gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n252), .A2(new_n254), .A3(new_n236), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n244), .B(new_n245), .C1(G183gat), .C2(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT25), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n219), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n219), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT25), .B1(new_n241), .B2(new_n247), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n255), .B1(new_n258), .B2(KEYINPUT25), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n265), .B2(new_n239), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n216), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n219), .ZN(new_n268));
  INV_X1    g067(.A(new_n216), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT29), .B1(new_n265), .B2(new_n239), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(new_n219), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT74), .B(new_n216), .C1(new_n262), .C2(new_n266), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  INV_X1    g075(.A(G64gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G92gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT30), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(new_n284), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(G127gat), .A2(G134gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  AND2_X1   g096(.A1(G127gat), .A2(G134gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G127gat), .A2(G134gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G113gat), .A2(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n296), .B(new_n300), .C1(new_n304), .C2(KEYINPUT1), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  AND2_X1   g106(.A1(G113gat), .A2(G120gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT68), .B1(new_n308), .B2(new_n301), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n295), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n305), .A2(new_n314), .A3(KEYINPUT80), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  OR2_X1    g119(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n319), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT79), .B(G162gat), .Z(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT2), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n322), .ZN(new_n330));
  NOR2_X1   g129(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n331));
  OAI21_X1  g130(.A(G141gat), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n324), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n326), .A2(new_n329), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n334), .A2(KEYINPUT76), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(G155gat), .B2(G162gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n336), .B(new_n337), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n317), .A2(new_n318), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n305), .A2(new_n314), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n343), .A2(new_n335), .A3(new_n341), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n293), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n345), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT83), .B1(new_n345), .B2(KEYINPUT5), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n335), .A2(new_n341), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(KEYINPUT81), .A3(new_n350), .A4(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n341), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT4), .B1(new_n352), .B2(new_n315), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n343), .A2(new_n335), .A3(new_n350), .A4(new_n341), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n317), .A2(new_n318), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n360), .A3(new_n341), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n292), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n357), .A2(new_n365), .A3(new_n292), .A4(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n348), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT0), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(G57gat), .ZN(new_n370));
  INV_X1    g169(.A(G85gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n354), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n362), .A3(new_n374), .A4(new_n292), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT84), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n372), .B1(new_n367), .B2(new_n376), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n367), .A2(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(new_n372), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n291), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT31), .B(G50gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G106gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n210), .A2(new_n215), .A3(new_n261), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT86), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n210), .A2(new_n215), .A3(new_n392), .A4(new_n261), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n360), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n352), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n361), .A2(new_n261), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n216), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G22gat), .B(G78gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n398), .B(KEYINPUT85), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n269), .B1(new_n361), .B2(new_n261), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n213), .A2(new_n211), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n261), .B1(new_n213), .B2(new_n211), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n360), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n352), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n400), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n402), .B1(new_n400), .B2(new_n409), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n389), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n401), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n400), .A2(new_n402), .A3(new_n409), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n388), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n382), .A2(new_n383), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n378), .A3(new_n377), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n275), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n260), .A2(new_n261), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n263), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n269), .B1(new_n424), .B2(new_n268), .ZN(new_n425));
  INV_X1    g224(.A(new_n271), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT37), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT87), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(KEYINPUT37), .C1(new_n425), .C2(new_n426), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n422), .A2(new_n428), .A3(new_n280), .A4(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT38), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n273), .A2(KEYINPUT37), .A3(new_n274), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n422), .A2(KEYINPUT38), .A3(new_n280), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n420), .A2(new_n436), .A3(new_n384), .A4(new_n282), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n292), .B1(new_n373), .B2(new_n362), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n342), .A2(new_n344), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n439), .B(KEYINPUT39), .C1(new_n293), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT39), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n383), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT40), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n445), .A2(new_n447), .B1(new_n382), .B2(new_n383), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n418), .B1(new_n448), .B2(new_n290), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n386), .A2(new_n418), .B1(new_n437), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G227gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n218), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n260), .A2(new_n343), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n315), .B1(new_n265), .B2(new_n239), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n260), .A2(new_n343), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n265), .A2(new_n315), .A3(new_n239), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(KEYINPUT32), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(G71gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(G99gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n459), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n471));
  INV_X1    g270(.A(new_n469), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(new_n462), .A3(new_n460), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n470), .B2(new_n473), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(KEYINPUT36), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT88), .B(new_n417), .C1(new_n474), .C2(new_n475), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n291), .C1(new_n381), .C2(new_n385), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n420), .A2(new_n384), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n291), .A4(new_n483), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n450), .A2(new_n481), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G127gat), .B(G155gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(G1gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT16), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G1gat), .B2(new_n491), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498));
  INV_X1    g297(.A(G57gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT93), .B1(new_n499), .B2(G64gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n277), .A3(G57gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(G64gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT9), .ZN(new_n506));
  NAND2_X1  g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n507), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n505), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT9), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n497), .B1(new_n498), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT96), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n517), .A2(new_n519), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n490), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  INV_X1    g323(.A(new_n490), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n515), .A2(new_n498), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G183gat), .B(G211gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT94), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT95), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n529), .B(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n523), .A2(new_n526), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n523), .B2(new_n526), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G190gat), .B(G218gat), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT98), .B1(new_n541), .B2(KEYINPUT7), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n546), .A2(new_n547), .A3(G85gat), .A4(G92gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(KEYINPUT97), .A3(KEYINPUT7), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n544), .A2(new_n545), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(G99gat), .B(G106gat), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n553), .B1(new_n371), .B2(new_n279), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n550), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT14), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n560), .B(new_n566), .C1(new_n562), .C2(new_n563), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n565), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n573), .A2(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n571), .B(new_n575), .C1(new_n570), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n560), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n558), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n584), .B(new_n585), .C1(new_n579), .C2(new_n558), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n537), .A2(new_n538), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT100), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n592), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n540), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n586), .A2(new_n587), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n591), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n539), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n536), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n489), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n551), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n509), .A2(new_n514), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n555), .B2(new_n556), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n550), .A2(new_n554), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n551), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n509), .A2(new_n514), .A3(new_n603), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT102), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n605), .A2(new_n610), .A3(new_n614), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n558), .A2(new_n611), .A3(new_n515), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n610), .ZN(new_n622));
  INV_X1    g421(.A(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT103), .Z(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(new_n251), .ZN(new_n627));
  INV_X1    g426(.A(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n621), .A2(KEYINPUT104), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n623), .B1(new_n616), .B2(new_n618), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n625), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n629), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(KEYINPUT105), .A3(new_n629), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n632), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n497), .B1(new_n582), .B2(new_n583), .ZN(new_n643));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n579), .ZN(new_n645));
  INV_X1    g444(.A(new_n497), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT92), .B1(new_n579), .B2(new_n497), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n644), .B(KEYINPUT13), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n645), .A2(KEYINPUT92), .A3(new_n646), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n643), .A2(KEYINPUT18), .A3(new_n644), .A4(new_n647), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n650), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G197gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT11), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n250), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT12), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n650), .A2(new_n663), .A3(new_n656), .A4(new_n657), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n642), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n601), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n486), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n492), .ZN(G1324gat));
  INV_X1    g471(.A(new_n670), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n290), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT16), .B(G8gat), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n674), .A2(KEYINPUT106), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(KEYINPUT106), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n675), .B1(new_n680), .B2(new_n676), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n680), .B2(G8gat), .ZN(new_n683));
  AOI211_X1 g482(.A(KEYINPUT107), .B(new_n496), .C1(new_n678), .C2(new_n679), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n677), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(G15gat), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n686), .A3(new_n481), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n673), .A2(new_n477), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n670), .A2(new_n417), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n595), .A2(new_n599), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n489), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n536), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n669), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n486), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n562), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n489), .B2(new_n694), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n386), .A2(new_n418), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n437), .A2(new_n449), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n481), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n485), .A2(new_n488), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n693), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n640), .A2(new_n641), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n631), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n667), .A3(new_n696), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT109), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n719), .B(new_n716), .C1(new_n702), .C2(new_n709), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n486), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n722), .ZN(G1328gat));
  NAND2_X1  g522(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n698), .A2(new_n563), .A3(new_n290), .A4(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n721), .B2(new_n291), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n708), .B1(new_n707), .B2(new_n693), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT44), .B(new_n694), .C1(new_n705), .C2(new_n706), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n717), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n719), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n710), .A2(KEYINPUT109), .A3(new_n717), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n481), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n730), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n698), .A2(new_n737), .A3(new_n477), .ZN(new_n739));
  INV_X1    g538(.A(new_n481), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n718), .B2(new_n720), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(KEYINPUT111), .A3(G43gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G43gat), .B1(new_n733), .B2(new_n481), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n739), .A3(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1330gat));
  OAI21_X1  g547(.A(G50gat), .B1(new_n733), .B2(new_n417), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n417), .A2(G50gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT112), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n698), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(KEYINPUT48), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n418), .B1(new_n718), .B2(new_n720), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n754), .A2(G50gat), .B1(new_n698), .B2(new_n751), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g555(.A(new_n715), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n600), .A2(new_n667), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(new_n707), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n699), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n290), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT113), .Z(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n759), .A2(new_n767), .A3(new_n477), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n759), .A2(new_n740), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n767), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g570(.A1(new_n759), .A2(new_n418), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n695), .A2(KEYINPUT115), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n667), .A2(new_n536), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n489), .B2(new_n694), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n775), .A4(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(new_n371), .A3(new_n699), .A4(new_n712), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n731), .A2(new_n732), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n775), .A2(new_n712), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT114), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n486), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n790), .ZN(G1336gat));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n290), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT116), .B1(new_n792), .B2(G92gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n715), .A2(G92gat), .A3(new_n291), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n782), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g596(.A1(new_n642), .A2(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n477), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n788), .A2(KEYINPUT117), .A3(new_n740), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n710), .A2(new_n740), .A3(new_n786), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(G99gat), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT118), .ZN(G1338gat));
  NOR2_X1   g605(.A1(new_n715), .A2(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n782), .A2(new_n418), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G106gat), .B1(new_n789), .B2(new_n417), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g610(.A1(new_n758), .A2(new_n642), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AOI211_X1 g612(.A(new_n620), .B(new_n617), .C1(new_n613), .C2(new_n615), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n634), .B1(new_n814), .B2(KEYINPUT119), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n616), .A2(new_n623), .A3(new_n618), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n630), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n635), .B1(new_n619), .B2(new_n620), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n617), .B1(new_n613), .B2(new_n615), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(KEYINPUT104), .A3(new_n623), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n813), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n817), .A2(new_n818), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(KEYINPUT119), .A3(new_n623), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n826), .A2(new_n621), .A3(KEYINPUT54), .A4(new_n827), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n813), .A2(new_n824), .A3(new_n629), .A4(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n631), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n644), .B1(new_n643), .B2(new_n647), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n654), .B1(new_n652), .B2(new_n655), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n662), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n666), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n694), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  INV_X1    g635(.A(new_n834), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n712), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n824), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT55), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n813), .A3(new_n824), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n632), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n667), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n642), .B2(new_n834), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n838), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n835), .B1(new_n845), .B2(new_n694), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n812), .B1(new_n846), .B2(new_n536), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n486), .A2(new_n290), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n476), .A2(new_n418), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n667), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(G113gat), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n851), .B2(new_n715), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n642), .A2(G120gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n851), .B2(new_n856), .ZN(G1341gat));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n536), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G127gat), .ZN(G1342gat));
  AOI211_X1 g658(.A(new_n694), .B(new_n851), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n830), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT121), .B(new_n631), .C1(new_n825), .C2(new_n829), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n667), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n712), .A2(new_n837), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n693), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n696), .B1(new_n869), .B2(new_n835), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n812), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n863), .B1(new_n871), .B2(new_n418), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n847), .A2(new_n863), .A3(new_n418), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n665), .A2(new_n666), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n481), .A2(new_n848), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n320), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n740), .A2(new_n417), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT122), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(KEYINPUT122), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n849), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n667), .A2(new_n320), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  OAI221_X1 g684(.A(new_n885), .B1(new_n881), .B2(new_n882), .C1(new_n876), .C2(new_n320), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1344gat));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n812), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n758), .A2(KEYINPUT123), .A3(new_n642), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n417), .B1(new_n870), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT124), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n847), .A2(KEYINPUT57), .A3(new_n418), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  INV_X1    g695(.A(new_n835), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n874), .B1(new_n830), .B2(new_n864), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n898), .A2(new_n866), .B1(new_n712), .B2(new_n837), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n899), .B2(new_n693), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(new_n696), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n895), .B(new_n863), .C1(new_n901), .C2(new_n417), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n893), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n712), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT59), .B(G148gat), .C1(new_n904), .C2(new_n875), .ZN(new_n905));
  INV_X1    g704(.A(new_n881), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n321), .A2(new_n322), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n712), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n909), .B2(new_n712), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n905), .B(new_n908), .C1(KEYINPUT59), .C2(new_n910), .ZN(G1345gat));
  AOI21_X1  g710(.A(G155gat), .B1(new_n906), .B2(new_n536), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n696), .A2(new_n328), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n909), .B2(new_n913), .ZN(G1346gat));
  NAND2_X1  g713(.A1(new_n906), .A2(new_n693), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n694), .A2(new_n327), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n915), .A2(new_n327), .B1(new_n909), .B2(new_n916), .ZN(G1347gat));
  AND2_X1   g716(.A1(new_n847), .A2(new_n486), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n290), .A3(new_n850), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(G169gat), .A3(new_n874), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  OAI21_X1  g720(.A(G169gat), .B1(new_n919), .B2(new_n874), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(new_n251), .B1(new_n919), .B2(new_n642), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n918), .A2(new_n850), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n715), .A2(new_n251), .A3(new_n291), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n927), .A2(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1349gat));
  OR3_X1    g730(.A1(new_n919), .A2(new_n696), .A3(new_n225), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n220), .B1(new_n919), .B2(new_n696), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1350gat));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G190gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n919), .A2(new_n694), .ZN(new_n940));
  MUX2_X1   g739(.A(new_n938), .B(new_n939), .S(new_n940), .Z(G1351gat));
  NOR3_X1   g740(.A1(new_n740), .A2(new_n699), .A3(new_n291), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n903), .A2(new_n667), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G197gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n918), .A2(new_n290), .A3(new_n878), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n874), .A2(G197gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  NOR3_X1   g746(.A1(new_n945), .A2(G204gat), .A3(new_n642), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n903), .A2(new_n757), .A3(new_n942), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n950), .B(new_n951), .C1(new_n628), .C2(new_n952), .ZN(G1353gat));
  OR3_X1    g752(.A1(new_n945), .A2(G211gat), .A3(new_n696), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n903), .A2(new_n536), .A3(new_n942), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1354gat));
  NAND4_X1  g757(.A1(new_n903), .A2(G218gat), .A3(new_n693), .A4(new_n942), .ZN(new_n959));
  INV_X1    g758(.A(G218gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n945), .B2(new_n694), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n959), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1355gat));
endmodule


