//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  NOR2_X1   g0015(.A1(new_n211), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n218), .B(new_n224), .C1(new_n213), .C2(new_n212), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n215), .A2(new_n225), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(G50), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(new_n221), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  MUX2_X1   g0048(.A(G226), .B(G232), .S(G1698), .Z(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n248), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT13), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n245), .B2(new_n246), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n258), .B(new_n259), .C1(new_n264), .C2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n268), .A3(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n268), .A3(G45), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G238), .A4(new_n247), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n255), .A2(new_n256), .A3(new_n265), .A4(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n249), .A2(new_n250), .B1(G33), .B2(G97), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n265), .B(new_n271), .C1(new_n273), .C2(new_n247), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT14), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT76), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(G179), .A3(new_n281), .A4(new_n272), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n276), .A2(new_n283), .A3(G169), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n221), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n222), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT71), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n222), .A2(KEYINPUT71), .A3(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n288), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n266), .A2(new_n268), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n287), .B1(new_n299), .B2(G20), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(KEYINPUT11), .B1(new_n300), .B2(G68), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n266), .A2(new_n268), .A3(G13), .A4(G20), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n301), .B(new_n305), .C1(KEYINPUT11), .C2(new_n297), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n285), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(G200), .B2(new_n276), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n280), .A2(G190), .A3(new_n281), .A4(new_n272), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(KEYINPUT73), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(KEYINPUT73), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n294), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G87), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT74), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(new_n324), .A3(new_n222), .A4(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G20), .A2(G77), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n317), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n287), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n302), .A2(G77), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n300), .B2(G77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n269), .A2(new_n270), .A3(new_n247), .ZN(new_n332));
  INV_X1    g0132(.A(G244), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n265), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n250), .A2(G238), .A3(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n250), .A2(G232), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G107), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(new_n250), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n248), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT72), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n265), .B(new_n342), .C1(new_n332), .C2(new_n333), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n331), .B1(G200), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n344), .A2(new_n348), .B1(new_n328), .B2(new_n330), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n335), .A2(new_n341), .A3(new_n343), .A4(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n345), .A2(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n313), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n314), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G58), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n302), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n358), .B2(new_n300), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT16), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT7), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G20), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n252), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G33), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT77), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n250), .B2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n356), .A2(new_n295), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n201), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n294), .A2(G159), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n295), .B1(new_n370), .B2(new_n371), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT78), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n362), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n367), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n222), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(new_n363), .B1(new_n385), .B2(new_n364), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT16), .B(new_n379), .C1(new_n387), .C2(new_n295), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n287), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n361), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n269), .A2(new_n270), .A3(G232), .A4(new_n247), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G223), .A2(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(G226), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(G1698), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n250), .B1(G33), .B2(G87), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n265), .B(new_n392), .C1(new_n396), .C2(new_n247), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(G190), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n397), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT17), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n397), .A2(new_n350), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(G169), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n391), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n380), .A2(new_n381), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n379), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n389), .B1(new_n413), .B2(new_n362), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n409), .B(new_n410), .C1(new_n414), .C2(new_n361), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n401), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n404), .A2(new_n408), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n300), .A2(G50), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G50), .B2(new_n302), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n355), .A2(new_n357), .A3(new_n291), .A4(new_n292), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n294), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n288), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G222), .A2(G1698), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n337), .A2(G223), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n250), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n248), .C1(G77), .C2(new_n250), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n265), .C1(new_n394), .C2(new_n332), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n346), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G200), .B2(new_n431), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n418), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n426), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n433), .ZN(new_n437));
  INV_X1    g0237(.A(new_n424), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n431), .A2(G179), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n431), .A2(new_n348), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n436), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n353), .A2(new_n417), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n302), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n266), .A2(new_n268), .A3(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n302), .A2(new_n288), .A3(new_n447), .A4(G116), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n286), .A2(new_n221), .B1(G20), .B2(new_n445), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(G33), .B2(G283), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G33), .B2(new_n253), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT20), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n446), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n384), .A2(new_n367), .A3(G264), .A4(G1698), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n384), .A2(new_n367), .A3(G257), .A4(new_n337), .ZN(new_n456));
  INV_X1    g0256(.A(G303), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(new_n456), .C1(new_n457), .C2(new_n250), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n248), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n266), .A2(new_n268), .A3(new_n460), .A4(G45), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n258), .ZN(new_n464));
  OAI211_X1 g0264(.A(G270), .B(new_n247), .C1(new_n461), .C2(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n454), .B1(new_n466), .B2(G200), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(KEYINPUT83), .B1(G190), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n454), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n468), .B2(new_n399), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n470), .A2(new_n466), .A3(new_n350), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n454), .A2(G169), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT21), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n466), .A2(new_n454), .A3(new_n478), .A4(G169), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n270), .A2(G250), .A3(new_n247), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n270), .A2(new_n247), .A3(KEYINPUT79), .A4(G250), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n333), .A2(G1698), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G238), .B2(G1698), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(new_n385), .ZN(new_n490));
  INV_X1    g0290(.A(new_n270), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n248), .B1(new_n491), .B2(new_n258), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(new_n492), .A3(G179), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n348), .B1(new_n486), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT80), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n486), .A2(new_n492), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G169), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT80), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n500));
  NAND3_X1  g0300(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n222), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n318), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n222), .A2(new_n501), .B1(new_n503), .B2(new_n318), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT81), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n384), .A2(new_n367), .A3(new_n222), .A4(G68), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n289), .B2(new_n253), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n321), .A2(new_n324), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(new_n287), .B1(new_n444), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  INV_X1    g0316(.A(new_n514), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n302), .A2(new_n288), .A3(new_n447), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT82), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n496), .A2(new_n500), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n486), .A2(G190), .A3(new_n492), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n399), .B1(new_n486), .B2(new_n492), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n519), .A2(G87), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n515), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n384), .A2(new_n367), .A3(new_n222), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n250), .A2(new_n532), .A3(new_n222), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n487), .A2(G20), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT84), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n222), .B2(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT23), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n537), .B(new_n540), .C1(new_n222), .C2(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n536), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n534), .A2(new_n535), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n535), .B1(new_n534), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n287), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n444), .A2(KEYINPUT25), .A3(new_n339), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT25), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n302), .B2(G107), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n548), .B1(new_n519), .B2(G107), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n384), .A2(new_n367), .A3(G257), .A4(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n384), .A2(new_n367), .A3(G250), .A4(new_n337), .ZN(new_n551));
  INV_X1    g0351(.A(G294), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n252), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n248), .ZN(new_n554));
  OAI211_X1 g0354(.A(G264), .B(new_n247), .C1(new_n461), .C2(new_n462), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n464), .A3(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n556), .A2(new_n399), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(G190), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n545), .B(new_n549), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n302), .A2(G97), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n253), .B2(new_n518), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n372), .A2(G107), .ZN(new_n563));
  XNOR2_X1  g0363(.A(G97), .B(G107), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n565), .A2(new_n253), .A3(G107), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n562), .B1(new_n571), .B2(new_n287), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n384), .A2(new_n367), .A3(G244), .A4(new_n337), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT4), .A2(G244), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1698), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n250), .A2(new_n578), .B1(G33), .B2(G283), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n248), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(new_n247), .C1(new_n461), .C2(new_n462), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n464), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(G190), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n580), .A2(new_n248), .B1(new_n258), .B2(new_n463), .ZN(new_n585));
  AOI21_X1  g0385(.A(G200), .B1(new_n585), .B2(new_n582), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(new_n348), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n294), .A2(G77), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n567), .B1(new_n565), .B2(new_n564), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(new_n222), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n339), .B1(new_n370), .B2(new_n371), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n287), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n562), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n585), .A2(new_n350), .A3(new_n582), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n559), .A2(new_n587), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n556), .A2(new_n348), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G179), .B2(new_n556), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n545), .B2(new_n549), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n443), .A2(new_n481), .A3(new_n529), .A4(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n498), .A2(new_n493), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n522), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n515), .B2(new_n527), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n510), .B(new_n512), .C1(new_n508), .C2(KEYINPUT81), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n505), .A2(new_n506), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n287), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n514), .A2(new_n444), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n607), .A2(new_n611), .A3(new_n612), .A4(new_n527), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n526), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(new_n559), .A3(new_n587), .A4(new_n597), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n545), .A2(new_n549), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n599), .C1(G179), .C2(new_n556), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n480), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n606), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n588), .A2(new_n595), .A3(new_n596), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n523), .A2(new_n528), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n614), .A2(new_n605), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT26), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(new_n621), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n443), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n441), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n408), .A2(new_n415), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n349), .A2(new_n351), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n308), .B1(new_n311), .B2(new_n632), .ZN(new_n633));
  NOR4_X1   g0433(.A1(new_n414), .A2(new_n400), .A3(new_n403), .A4(new_n361), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT17), .B1(new_n391), .B2(new_n401), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n630), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n436), .A2(new_n437), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n628), .A2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(G330), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n222), .A2(G13), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n299), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT86), .B1(new_n644), .B2(KEYINPUT27), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT86), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT27), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n299), .A2(new_n646), .A3(new_n647), .A4(new_n643), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G213), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n644), .B2(KEYINPUT27), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n649), .A2(G343), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n481), .B1(new_n470), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n477), .A2(new_n479), .ZN(new_n655));
  INV_X1    g0455(.A(new_n475), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n454), .A3(new_n652), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n642), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n601), .A2(new_n653), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n617), .A2(new_n652), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n559), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n662), .B2(new_n601), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n480), .A2(new_n652), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n664), .A2(new_n666), .B1(new_n601), .B2(new_n653), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n216), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n264), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n259), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n504), .A2(G116), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n670), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n219), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n675), .B2(KEYINPUT87), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(KEYINPUT87), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT89), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n622), .A2(new_n625), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n614), .A2(new_n621), .A3(KEYINPUT26), .A4(new_n605), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n620), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n683), .B2(new_n653), .ZN(new_n684));
  AOI211_X1 g0484(.A(KEYINPUT89), .B(new_n652), .C1(new_n620), .C2(new_n682), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT29), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n627), .A2(new_n653), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n602), .A2(new_n481), .A3(new_n529), .A4(new_n653), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n493), .A2(new_n466), .ZN(new_n692));
  INV_X1    g0492(.A(new_n583), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n554), .A2(new_n555), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT88), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n697), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n692), .A2(new_n693), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(G179), .B1(new_n486), .B2(new_n492), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n583), .A3(new_n466), .A4(new_n556), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n703), .B2(new_n652), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n691), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n690), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n678), .B1(new_n710), .B2(G1), .ZN(G364));
  INV_X1    g0511(.A(new_n659), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n654), .A2(new_n642), .A3(new_n658), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n643), .A2(G45), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n671), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT91), .Z(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n654), .A2(new_n658), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n717), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n250), .A2(new_n216), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n724), .A2(new_n725), .B1(G116), .B2(new_n216), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n243), .A2(G45), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n669), .A2(new_n250), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G45), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n220), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n726), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n221), .B1(G20), .B2(new_n348), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n721), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n723), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n737));
  NAND2_X1  g0537(.A1(G20), .A2(G179), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT93), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n399), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n346), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  AOI22_X1  g0543(.A1(G50), .A2(new_n741), .B1(new_n743), .B2(G77), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n740), .A2(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n742), .A2(new_n399), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n744), .B1(new_n356), .B2(new_n746), .C1(new_n295), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n222), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n346), .A3(new_n399), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n346), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n222), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n750), .A2(new_n346), .A3(G200), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n754), .B1(new_n253), .B2(new_n756), .C1(new_n339), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n318), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n749), .A2(new_n385), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G311), .A2(new_n743), .B1(new_n741), .B2(G326), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n748), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n756), .ZN(new_n765));
  INV_X1    g0565(.A(new_n751), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n765), .A2(G294), .B1(new_n766), .B2(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n767), .B1(new_n768), .B2(new_n757), .C1(new_n746), .C2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n385), .B1(new_n759), .B2(new_n457), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT94), .Z(new_n772));
  NOR3_X1   g0572(.A1(new_n764), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n733), .B1(new_n761), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n722), .A2(new_n737), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n718), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(G396));
  NAND2_X1  g0578(.A1(new_n331), .A2(new_n652), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n344), .A2(new_n348), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n780), .A2(new_n331), .A3(new_n652), .A4(new_n351), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT97), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n349), .A2(KEYINPUT97), .A3(new_n351), .A4(new_n652), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n352), .A2(new_n779), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n687), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n785), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n626), .A2(new_n623), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n657), .A2(new_n601), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n605), .B1(new_n789), .B2(new_n615), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n787), .B(new_n653), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n723), .B1(new_n792), .B2(new_n708), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n708), .B2(new_n792), .ZN(new_n794));
  INV_X1    g0594(.A(G77), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n733), .A2(new_n719), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n717), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G283), .A2(new_n747), .B1(new_n745), .B2(G294), .ZN(new_n798));
  INV_X1    g0598(.A(new_n741), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n457), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n385), .B1(new_n759), .B2(new_n339), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT95), .Z(new_n802));
  INV_X1    g0602(.A(new_n743), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n445), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n765), .A2(G97), .B1(new_n766), .B2(G311), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n318), .B2(new_n757), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n800), .A2(new_n802), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G143), .A2(new_n745), .B1(new_n743), .B2(G159), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G137), .A2(new_n741), .B1(new_n747), .B2(G150), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n250), .B1(new_n751), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT96), .Z(new_n814));
  OR2_X1    g0614(.A1(new_n757), .A2(new_n295), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n815), .B1(new_n202), .B2(new_n759), .C1(new_n356), .C2(new_n756), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n807), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n733), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n797), .B1(new_n818), .B2(new_n819), .C1(new_n787), .C2(new_n720), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n794), .A2(new_n820), .ZN(G384));
  OR2_X1    g0621(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(G116), .A3(new_n223), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  OAI21_X1  g0625(.A(G77), .B1(new_n356), .B2(new_n295), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n826), .A2(new_n219), .B1(G50), .B2(new_n295), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n299), .A2(G13), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n410), .B1(new_n414), .B2(new_n361), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n649), .A2(new_n651), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n414), .B2(new_n361), .ZN(new_n835));
  AND4_X1   g0635(.A1(new_n831), .A2(new_n832), .A3(new_n835), .A4(new_n402), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n407), .A2(new_n833), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n385), .A2(new_n364), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n371), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G68), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n840), .B2(new_n379), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n360), .B1(new_n389), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT98), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT98), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n844), .B(new_n360), .C1(new_n389), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n837), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n831), .B1(new_n846), .B2(new_n402), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n843), .A2(new_n845), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n834), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n630), .B2(new_n636), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n830), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n417), .A2(new_n834), .A3(new_n849), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n832), .A2(new_n835), .A3(new_n402), .A4(new_n831), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n846), .A2(new_n402), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n831), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n856), .A3(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n652), .A2(new_n306), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n307), .A2(new_n311), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n306), .B(new_n652), .C1(new_n312), .C2(new_n285), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n785), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n707), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n707), .A2(new_n862), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n832), .A2(new_n835), .A3(new_n402), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(new_n854), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n835), .B1(new_n630), .B2(new_n636), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n830), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n866), .B1(new_n871), .B2(new_n857), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n865), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n873), .A2(new_n443), .A3(new_n707), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n443), .B2(new_n707), .ZN(new_n875));
  OR3_X1    g0675(.A1(new_n874), .A2(new_n875), .A3(new_n642), .ZN(new_n876));
  INV_X1    g0676(.A(new_n835), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n417), .A2(new_n877), .B1(new_n868), .B2(new_n854), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n857), .B1(KEYINPUT38), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n307), .A2(new_n652), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n852), .A2(KEYINPUT39), .A3(new_n857), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n630), .A2(new_n834), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n860), .A2(new_n861), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n631), .A2(new_n652), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n791), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n885), .B1(new_n890), .B2(new_n858), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n686), .A2(new_n443), .A3(new_n689), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n640), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n892), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n876), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n299), .B2(new_n643), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n876), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n829), .B1(new_n897), .B2(new_n898), .ZN(G367));
  OAI211_X1 g0699(.A(new_n587), .B(new_n597), .C1(new_n572), .C2(new_n653), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n621), .A2(new_n652), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n902), .B(KEYINPUT99), .Z(new_n903));
  NOR2_X1   g0703(.A1(new_n665), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT100), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n608), .A2(new_n613), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n652), .ZN(new_n907));
  MUX2_X1   g0707(.A(new_n606), .B(new_n624), .S(new_n907), .Z(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n905), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n666), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n663), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n902), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT42), .Z(new_n914));
  OAI21_X1  g0714(.A(new_n597), .B1(new_n903), .B2(new_n618), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n653), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n914), .A2(new_n916), .B1(KEYINPUT43), .B2(new_n908), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n910), .A2(new_n917), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n920));
  XNOR2_X1  g0720(.A(new_n670), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n663), .A2(new_n911), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT102), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n659), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n659), .A2(new_n924), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n926), .A2(new_n927), .B1(new_n663), .B2(new_n911), .ZN(new_n928));
  INV_X1    g0728(.A(new_n927), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n912), .A3(new_n925), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n710), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n931), .A2(new_n708), .A3(new_n690), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT45), .ZN(new_n935));
  INV_X1    g0735(.A(new_n667), .ZN(new_n936));
  INV_X1    g0736(.A(new_n902), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n902), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(KEYINPUT44), .A3(new_n937), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT44), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n667), .B2(new_n902), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n665), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n940), .A2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(new_n665), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n932), .A2(new_n934), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n921), .B1(new_n949), .B2(new_n710), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n716), .A2(G1), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT104), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n918), .B(new_n919), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n230), .A2(new_n729), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n734), .B1(new_n216), .B2(new_n514), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n723), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n757), .A2(new_n795), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n385), .B(new_n957), .C1(G137), .C2(new_n766), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n756), .A2(new_n295), .ZN(new_n959));
  INV_X1    g0759(.A(new_n759), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(G58), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n747), .A2(G159), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n741), .A2(G143), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G50), .A2(new_n743), .B1(new_n745), .B2(G150), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G303), .A2(new_n745), .B1(new_n741), .B2(G311), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n757), .A2(new_n253), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n385), .B1(new_n751), .B2(new_n970), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(G107), .C2(new_n765), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n960), .A2(G116), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT46), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G283), .A2(new_n743), .B1(new_n747), .B2(G294), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n968), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n966), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n956), .B1(new_n979), .B2(new_n733), .ZN(new_n980));
  INV_X1    g0780(.A(new_n721), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n908), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n953), .A2(new_n982), .ZN(G387));
  NAND2_X1  g0783(.A1(new_n932), .A2(new_n934), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n670), .C1(new_n710), .C2(new_n931), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n315), .A2(new_n316), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n202), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(G45), .B1(G68), .B2(G77), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n672), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n988), .B1(new_n987), .B2(new_n202), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n728), .B1(new_n730), .B2(new_n234), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(G107), .B2(new_n216), .C1(new_n672), .C2(new_n724), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n717), .B1(new_n994), .B2(new_n734), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n664), .B2(new_n981), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n385), .B(new_n969), .C1(G150), .C2(new_n766), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n517), .A2(new_n765), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n960), .A2(G77), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n202), .A2(new_n746), .B1(new_n799), .B2(new_n752), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n358), .A2(new_n748), .B1(new_n803), .B2(new_n295), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n250), .B1(new_n766), .B2(G326), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n756), .A2(new_n768), .B1(new_n759), .B2(new_n552), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G311), .A2(new_n747), .B1(new_n741), .B2(G322), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n457), .B2(new_n803), .C1(new_n970), .C2(new_n746), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT48), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT49), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1005), .B1(new_n445), .B2(new_n757), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1004), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n996), .B1(new_n1015), .B2(new_n733), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n952), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n928), .B2(new_n930), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT106), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT106), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n985), .A2(new_n1021), .ZN(G393));
  AOI21_X1  g0822(.A(new_n735), .B1(G97), .B2(new_n669), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n239), .A2(new_n728), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n717), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G311), .A2(new_n745), .B1(new_n741), .B2(G317), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT52), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n756), .A2(new_n445), .B1(new_n759), .B2(new_n768), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n385), .B1(new_n751), .B2(new_n769), .C1(new_n339), .C2(new_n757), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G303), .C2(new_n747), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n552), .B2(new_n803), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n385), .B1(new_n766), .B2(G143), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n318), .B2(new_n757), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G150), .A2(new_n741), .B1(new_n745), .B2(G159), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT51), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1034), .B(new_n1036), .C1(G68), .C2(new_n960), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n756), .A2(new_n795), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n748), .B2(new_n202), .C1(new_n986), .C2(new_n803), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT110), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1032), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1025), .B1(new_n1042), .B2(new_n819), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n903), .B2(new_n721), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n665), .B1(new_n940), .B2(new_n944), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1047), .B2(new_n952), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1045), .B(new_n948), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1049), .A2(new_n984), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n949), .A2(new_n670), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(G390));
  AND4_X1   g0852(.A1(KEYINPUT26), .A2(new_n614), .A3(new_n621), .A4(new_n605), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n625), .B2(new_n622), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n653), .B1(new_n1054), .B2(new_n790), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(KEYINPUT89), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n683), .A2(new_n679), .A3(new_n653), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n785), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT111), .B1(new_n1058), .B2(new_n888), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n787), .B1(new_n684), .B2(new_n685), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n889), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n886), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n882), .B1(new_n871), .B2(new_n857), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n706), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n704), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n642), .B1(new_n1067), .B2(new_n691), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1068), .A2(new_n787), .A3(new_n886), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT112), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(KEYINPUT112), .A3(new_n787), .A4(new_n886), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n890), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n882), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n881), .A2(new_n883), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1065), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n787), .B1(new_n1068), .B2(KEYINPUT113), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n707), .A2(KEYINPUT113), .A3(G330), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n887), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT114), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(KEYINPUT114), .B(new_n887), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1081), .A2(new_n1086), .A3(new_n1073), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n791), .A2(new_n889), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1069), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n886), .B1(new_n1068), .B2(new_n787), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n443), .A2(new_n1068), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n893), .A2(new_n640), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1080), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n1078), .C1(new_n1069), .C2(new_n1079), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1100), .A3(new_n670), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1078), .B(new_n952), .C1(new_n1069), .C2(new_n1079), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n250), .B(new_n760), .C1(G294), .C2(new_n766), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n815), .A3(new_n1039), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G97), .A2(new_n743), .B1(new_n741), .B2(G283), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n339), .B2(new_n748), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G116), .C2(new_n745), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n960), .A2(G150), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT53), .Z(new_n1111));
  AOI22_X1  g0911(.A1(G128), .A2(new_n741), .B1(new_n747), .B2(G137), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT54), .B(G143), .Z(new_n1113));
  AOI22_X1  g0913(.A1(G132), .A2(new_n745), .B1(new_n743), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n250), .B1(new_n751), .B2(new_n1115), .C1(new_n202), .C2(new_n757), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G159), .B2(new_n765), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1109), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n733), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n717), .B1(new_n358), .B2(new_n796), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT115), .Z(new_n1123));
  AND2_X1   g0923(.A1(new_n881), .A2(new_n883), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1123), .C1(new_n1124), .C2(new_n720), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1102), .A2(KEYINPUT117), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT117), .B1(new_n1102), .B2(new_n1125), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1101), .B1(new_n1126), .B2(new_n1127), .ZN(G378));
  NOR2_X1   g0928(.A1(new_n424), .A2(new_n833), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n639), .A2(new_n441), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n442), .A2(new_n1129), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n866), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n863), .B1(new_n879), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n707), .A2(new_n862), .A3(new_n863), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n857), .B2(new_n852), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1138), .B(G330), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1138), .B1(new_n873), .B2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n892), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(G330), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1138), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n884), .A2(new_n891), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1143), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1151), .A3(KEYINPUT122), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT122), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n892), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1138), .A2(new_n720), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n765), .A2(G150), .B1(new_n960), .B2(new_n1113), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n748), .B2(new_n812), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n745), .A2(G128), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n799), .B2(new_n1115), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G137), .C2(new_n743), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT120), .Z(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  AOI211_X1 g0964(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n752), .B2(new_n757), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n264), .A2(new_n250), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n959), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n766), .A2(G283), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1171), .A2(new_n999), .A3(new_n1168), .A4(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G116), .A2(new_n741), .B1(new_n743), .B2(new_n517), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n757), .A2(new_n356), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT118), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(new_n339), .C2(new_n746), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1173), .B(new_n1177), .C1(G97), .C2(new_n747), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1170), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1180), .B2(new_n1178), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n733), .B1(new_n1167), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT121), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n717), .B1(new_n202), .B2(new_n796), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1155), .A2(new_n952), .B1(new_n1156), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1069), .B1(new_n1065), .B2(new_n1077), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1189), .B(new_n1076), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1095), .B1(new_n1191), .B2(new_n1099), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT123), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1146), .A2(new_n1151), .A3(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT123), .A4(new_n1143), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n670), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1096), .B1(new_n1080), .B2(new_n1097), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1198), .B2(new_n1155), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1187), .B1(new_n1197), .B2(new_n1199), .ZN(G375));
  INV_X1    g1000(.A(new_n921), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1097), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n887), .A2(new_n719), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n733), .A2(G68), .A3(new_n719), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G283), .A2(new_n745), .B1(new_n741), .B2(G294), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G107), .A2(new_n743), .B1(new_n747), .B2(G116), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n385), .B1(new_n751), .B2(new_n457), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n957), .B(new_n1208), .C1(G97), .C2(new_n960), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n998), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1176), .A2(new_n250), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT124), .Z(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n766), .B1(new_n960), .B2(G159), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n202), .B2(new_n756), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n747), .B2(new_n1113), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G137), .A2(new_n745), .B1(new_n743), .B2(G150), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n812), .C2(new_n799), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n717), .B(new_n1205), .C1(new_n1218), .C2(new_n733), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1093), .A2(new_n952), .B1(new_n1204), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1203), .A2(new_n1220), .ZN(G381));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G393), .A2(G396), .ZN(new_n1223));
  INV_X1    g1023(.A(G384), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G387), .A3(G381), .ZN(new_n1226));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1102), .A2(new_n1125), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n674), .B1(new_n1080), .B2(new_n1097), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n1100), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(G407));
  NOR2_X1   g1031(.A1(new_n650), .A2(G343), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT125), .Z(new_n1233));
  NAND3_X1  g1033(.A1(new_n1227), .A2(new_n1230), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1095), .A4(new_n1092), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n670), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1239), .B2(new_n1202), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1220), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1224), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1202), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(KEYINPUT60), .B2(new_n1097), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1220), .B(G384), .C1(new_n1244), .C2(new_n1238), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G378), .B(new_n1187), .C1(new_n1199), .C2(new_n1197), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1198), .A2(new_n1201), .A3(new_n1155), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1194), .A2(new_n952), .A3(new_n1195), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1186), .A2(new_n1156), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1230), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1232), .B(new_n1246), .C1(new_n1247), .C2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1236), .B1(new_n1253), .B2(KEYINPUT63), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n777), .B1(new_n985), .B2(new_n1021), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1223), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n953), .A2(G390), .A3(new_n982), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G390), .B1(new_n953), .B2(new_n982), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1222), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1233), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1246), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G378), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1252), .B1(G375), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1232), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1246), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(KEYINPUT126), .A3(new_n1267), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1242), .A2(new_n1245), .B1(G2897), .B2(new_n1233), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1232), .A2(G2897), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1246), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1254), .A2(new_n1269), .A3(new_n1275), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1246), .A2(new_n1283), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1274), .A2(new_n1283), .B1(new_n1266), .B2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1279), .A2(new_n1277), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1262), .B1(new_n1286), .B2(new_n1266), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1281), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1230), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1282), .A2(KEYINPUT127), .A3(new_n1246), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1227), .A2(G378), .B1(new_n1273), .B2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1261), .B(new_n1264), .C1(new_n1292), .C2(new_n1273), .ZN(new_n1294));
  AND4_X1   g1094(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1291), .A2(new_n1294), .B1(new_n1293), .B2(new_n1290), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


