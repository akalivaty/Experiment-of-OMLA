//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT70), .B1(new_n189), .B2(G116), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(new_n187), .A3(G119), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  AND2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n193), .A2(new_n194), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT0), .B(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(KEYINPUT0), .A3(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n201), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT71), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n214), .B2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n216), .A2(new_n222), .A3(new_n218), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n201), .A2(new_n210), .A3(new_n225), .A4(new_n211), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n213), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  AOI21_X1  g042(.A(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n204), .A2(KEYINPUT1), .A3(G146), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n228), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT67), .B(new_n230), .C1(new_n199), .C2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n206), .A2(KEYINPUT1), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n219), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n239), .B2(new_n215), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n227), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n198), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(KEYINPUT68), .A3(new_n242), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n236), .B1(new_n232), .B2(new_n233), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(new_n241), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n212), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n201), .A2(new_n210), .A3(KEYINPUT65), .A4(new_n211), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n224), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n253), .A2(new_n224), .A3(new_n257), .A4(new_n254), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n245), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n245), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n246), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n227), .A2(new_n243), .A3(new_n197), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT72), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n227), .A2(new_n243), .A3(new_n267), .A4(new_n197), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n270), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n274), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n264), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n246), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n245), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n259), .B2(new_n245), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n278), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n250), .A2(new_n247), .B1(new_n255), .B2(KEYINPUT66), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n197), .B1(new_n288), .B2(new_n258), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n266), .A2(new_n268), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT28), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n277), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n262), .A2(new_n263), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n278), .B1(new_n295), .B2(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT32), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n291), .A2(new_n277), .A3(new_n293), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n277), .B1(new_n283), .B2(new_n269), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n244), .A2(new_n198), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n269), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT28), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n293), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n276), .A2(new_n306), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n276), .B1(new_n264), .B2(new_n290), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n306), .A4(new_n305), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n309), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  INV_X1    g133(.A(new_n300), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n287), .B2(new_n298), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT32), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n303), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  INV_X1    g139(.A(G902), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(G234), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n335), .B2(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(KEYINPUT78), .A3(new_n202), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n334), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G119), .B(G128), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT76), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT77), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n189), .B2(G128), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n349), .B(new_n350), .C1(G119), .C2(new_n235), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(G110), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT77), .B1(new_n345), .B2(new_n346), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n336), .A2(G146), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n337), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(G110), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n356), .B(new_n357), .C1(new_n345), .C2(new_n346), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n360), .B(new_n361), .Z(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT79), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n354), .A2(new_n358), .A3(new_n362), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT81), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT81), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n329), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n327), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(new_n326), .A3(new_n367), .ZN(new_n374));
  NOR2_X1   g188(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n375), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n365), .A2(new_n326), .A3(new_n367), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n324), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n371), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n328), .B1(new_n381), .B2(new_n369), .ZN(new_n382));
  INV_X1    g196(.A(new_n379), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT82), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n235), .A2(G143), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n204), .A2(G128), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n386), .A2(new_n387), .A3(G134), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n187), .A2(G122), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n204), .A2(G128), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n387), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(KEYINPUT13), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n214), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT96), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT97), .B1(new_n391), .B2(KEYINPUT14), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n390), .A3(new_n403), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n391), .A2(KEYINPUT97), .A3(KEYINPUT14), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G134), .B1(new_n386), .B2(new_n387), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n393), .B1(new_n388), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n400), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n393), .A2(new_n394), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n388), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n415), .A2(new_n325), .A3(G953), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n410), .A2(KEYINPUT98), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n401), .A3(new_n409), .ZN(new_n419));
  INV_X1    g233(.A(new_n416), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n326), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT99), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G478), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(KEYINPUT15), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(KEYINPUT99), .A3(new_n326), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n424), .B2(new_n428), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n204), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n432), .B(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n222), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(KEYINPUT17), .A3(G131), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n438), .A2(new_n355), .A3(new_n337), .A4(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT94), .B(G104), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g257(.A1(KEYINPUT18), .A2(G131), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n433), .B(new_n444), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n340), .A2(KEYINPUT92), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n340), .A2(KEYINPUT92), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G146), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n342), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(KEYINPUT19), .A3(new_n447), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n453), .B(new_n202), .C1(KEYINPUT19), .C2(new_n340), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n434), .A2(new_n436), .B1(G146), .B2(new_n336), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n450), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n443), .B1(new_n457), .B2(KEYINPUT93), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n454), .A2(new_n455), .B1(new_n445), .B2(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT93), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n452), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(G475), .A2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT20), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n461), .ZN(new_n466));
  INV_X1    g280(.A(new_n443), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n451), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n443), .B1(new_n440), .B2(new_n450), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n326), .B1(new_n452), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT95), .B(new_n326), .C1(new_n452), .C2(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(G475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n272), .A2(G952), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(G234), .B2(G237), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n326), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n431), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G210), .B1(G237), .B2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT8), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G104), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT85), .B1(new_n491), .B2(G107), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(G107), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n491), .A2(KEYINPUT85), .A3(G107), .ZN(new_n495));
  OAI21_X1  g309(.A(G101), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT3), .B1(new_n491), .B2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n392), .A3(G104), .ZN(new_n499));
  INV_X1    g313(.A(G101), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n493), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n189), .A2(G116), .ZN(new_n503));
  OAI21_X1  g317(.A(G113), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n193), .B2(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n195), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n502), .A2(new_n195), .A3(new_n505), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(KEYINPUT90), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n490), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n249), .A2(new_n333), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n212), .A2(G125), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT89), .B(G224), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n272), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n497), .A2(new_n499), .A3(new_n493), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n524), .A2(new_n526), .B1(new_n195), .B2(new_n196), .ZN(new_n527));
  INV_X1    g341(.A(new_n502), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n193), .A2(new_n194), .ZN(new_n529));
  INV_X1    g343(.A(new_n505), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n531), .A3(new_n488), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n513), .A2(KEYINPUT7), .A3(new_n514), .A4(new_n517), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n519), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n326), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n488), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n520), .A2(new_n523), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n193), .A2(new_n194), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n537), .A2(new_n525), .B1(new_n538), .B2(new_n529), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n508), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n540), .A3(KEYINPUT6), .ZN(new_n541));
  INV_X1    g355(.A(new_n517), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n515), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(new_n536), .C1(new_n539), .C2(new_n508), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n487), .B1(new_n535), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n519), .A2(new_n532), .A3(new_n533), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT90), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n506), .B1(new_n531), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n489), .B1(new_n552), .B2(new_n510), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n486), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(KEYINPUT91), .B2(new_n549), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n238), .A2(new_n528), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n230), .B1(new_n199), .B2(G128), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n236), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT86), .B(new_n230), .C1(new_n199), .C2(G128), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n502), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n224), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT12), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT87), .B(KEYINPUT10), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n565), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n237), .A2(new_n573), .A3(new_n568), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n574), .B2(new_n502), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n213), .B(new_n226), .C1(new_n524), .C2(new_n526), .ZN(new_n576));
  INV_X1    g390(.A(new_n224), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n238), .A2(KEYINPUT10), .A3(new_n528), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n224), .C1(new_n564), .C2(new_n569), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n272), .A2(G227), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT83), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n224), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n579), .A3(new_n586), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G469), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT88), .B(G469), .Z(new_n595));
  NOR2_X1   g409(.A1(new_n582), .A2(new_n587), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n586), .B1(new_n590), .B2(new_n579), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n326), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n563), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n485), .A2(new_n561), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n323), .A2(new_n385), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT100), .B(G101), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G3));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n299), .B2(new_n326), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n380), .A2(new_n599), .A3(new_n384), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n605), .A2(new_n606), .A3(new_n321), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n549), .A2(new_n556), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT101), .B1(new_n608), .B2(new_n559), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n610), .B(new_n560), .C1(new_n549), .C2(new_n556), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n484), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n416), .B(KEYINPUT102), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n419), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT103), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n617), .B(KEYINPUT33), .C1(new_n419), .C2(new_n420), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n423), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n618), .A2(G478), .A3(new_n326), .A4(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n479), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n607), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT105), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  INV_X1    g444(.A(new_n479), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n431), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n614), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n607), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT106), .B(KEYINPUT35), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NOR2_X1   g451(.A1(new_n605), .A2(new_n321), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n359), .B(KEYINPUT107), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n328), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n383), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n561), .A2(new_n485), .A3(new_n599), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  NAND3_X1  g462(.A1(new_n612), .A2(new_n599), .A3(new_n644), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n481), .B1(new_n482), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n649), .A2(new_n632), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n323), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  AOI21_X1  g468(.A(new_n604), .B1(new_n311), .B2(new_n276), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n279), .A2(new_n286), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(G472), .A2(G902), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n656), .A2(KEYINPUT108), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT108), .B1(new_n656), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n303), .A3(new_n322), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n651), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n599), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n431), .A2(new_n479), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n383), .A3(new_n559), .A4(new_n643), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n558), .B(KEYINPUT38), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n661), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  INV_X1    g485(.A(new_n651), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n623), .A2(new_n479), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n649), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n323), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  INV_X1    g490(.A(new_n596), .ZN(new_n677));
  INV_X1    g491(.A(new_n597), .ZN(new_n678));
  AOI21_X1  g492(.A(G902), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n598), .B(new_n562), .C1(new_n679), .C2(new_n593), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n323), .A2(new_n625), .A3(new_n385), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n323), .A2(new_n633), .A3(new_n385), .A4(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n535), .A2(new_n548), .A3(new_n487), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n486), .B1(new_n554), .B2(new_n555), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n559), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n610), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n608), .A2(KEYINPUT101), .A3(new_n559), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n687), .B1(new_n693), .B2(new_n680), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n612), .A2(new_n681), .A3(KEYINPUT109), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n323), .A2(new_n485), .A3(new_n644), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NAND2_X1  g512(.A1(new_n612), .A2(new_n665), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n699), .A2(new_n484), .A3(new_n680), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n372), .A2(new_n379), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n277), .B1(new_n312), .B2(new_n293), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n296), .B2(new_n297), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n320), .B1(new_n703), .B2(new_n287), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n299), .A2(new_n326), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT110), .B(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n700), .A2(new_n701), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  INV_X1    g523(.A(new_n673), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n696), .A2(new_n707), .A3(new_n644), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  NAND2_X1  g526(.A1(new_n588), .A2(new_n591), .ZN(new_n713));
  MUX2_X1   g527(.A(new_n713), .B(new_n591), .S(KEYINPUT111), .Z(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n593), .ZN(new_n715));
  INV_X1    g529(.A(new_n598), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n593), .A2(new_n326), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n558), .A2(new_n559), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n718), .A2(new_n563), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n323), .A2(new_n720), .A3(new_n385), .A4(new_n710), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n701), .ZN(new_n725));
  INV_X1    g539(.A(new_n319), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n299), .B2(new_n300), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n302), .B(new_n320), .C1(new_n287), .C2(new_n298), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT112), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n321), .B2(KEYINPUT32), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n726), .B1(new_n732), .B2(KEYINPUT113), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n734), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n725), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n710), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n724), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n222), .ZN(G33));
  NOR2_X1   g553(.A1(new_n632), .A2(new_n651), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n323), .A2(new_n720), .A3(new_n385), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n714), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n588), .B2(new_n591), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n593), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n717), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n598), .B1(new_n747), .B2(KEYINPUT46), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n562), .B(new_n662), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n479), .B1(new_n622), .B2(new_n621), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT43), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(new_n644), .C1(new_n321), .C2(new_n605), .ZN(new_n754));
  AOI211_X1 g568(.A(new_n719), .B(new_n750), .C1(new_n751), .C2(new_n754), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  OAI21_X1  g572(.A(new_n562), .B1(new_n748), .B2(new_n749), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT47), .Z(new_n760));
  NAND3_X1  g574(.A1(new_n558), .A2(new_n559), .A3(new_n672), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n323), .A2(new_n385), .A3(new_n624), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NAND2_X1  g578(.A1(new_n753), .A2(new_n481), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n680), .A3(new_n719), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n736), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n385), .A2(new_n481), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n661), .A2(new_n680), .A3(new_n769), .A4(new_n719), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n479), .A3(new_n623), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n707), .A2(new_n701), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n696), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(G952), .A3(new_n774), .A4(new_n272), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT121), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n759), .B(KEYINPUT47), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n598), .B1(new_n679), .B2(new_n593), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n563), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n765), .A2(new_n772), .A3(new_n719), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n668), .A2(new_n559), .A3(new_n680), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT50), .Z(new_n787));
  NOR2_X1   g601(.A1(new_n623), .A2(new_n479), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n707), .A2(new_n644), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n770), .A2(new_n788), .B1(new_n766), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n776), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n781), .B(KEYINPUT119), .Z(new_n793));
  NAND2_X1  g607(.A1(new_n778), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n783), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT120), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT120), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n791), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n768), .B(new_n792), .C1(new_n798), .C2(KEYINPUT51), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n682), .A2(new_n685), .A3(new_n697), .A4(new_n708), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n599), .A2(new_n644), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n801), .A2(new_n761), .A3(new_n431), .A4(new_n479), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n323), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n720), .A2(new_n644), .A3(new_n710), .A4(new_n707), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n741), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n632), .A2(new_n624), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n561), .A3(new_n613), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n607), .A2(new_n807), .B1(new_n638), .B2(new_n645), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n601), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n808), .B2(new_n601), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n800), .B(new_n805), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n738), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n323), .B1(new_n652), .B2(new_n674), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n563), .B1(new_n672), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n816), .B2(new_n672), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n644), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n718), .A2(new_n699), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n661), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n815), .A2(new_n821), .A3(new_n711), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n815), .A2(new_n821), .A3(KEYINPUT52), .A4(new_n711), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n828), .A3(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n814), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n832), .A3(new_n825), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n825), .A2(new_n832), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n814), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n733), .A2(new_n735), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n701), .A3(new_n737), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n723), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n682), .A2(new_n685), .A3(new_n697), .A4(new_n708), .ZN(new_n843));
  INV_X1    g657(.A(new_n812), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n810), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n845), .A3(new_n805), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n833), .A2(new_n834), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n837), .B(new_n839), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT54), .B1(new_n838), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n814), .A2(new_n835), .A3(KEYINPUT53), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n814), .A2(new_n830), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n799), .A2(new_n855), .B1(G952), .B2(G953), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n779), .B(KEYINPUT49), .Z(new_n857));
  NOR3_X1   g671(.A1(new_n725), .A2(new_n560), .A3(new_n563), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n752), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n859), .A2(new_n668), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n856), .B1(new_n661), .B2(new_n860), .ZN(G75));
  NOR2_X1   g675(.A1(new_n272), .A2(G952), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n852), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n814), .B2(new_n830), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n326), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n867), .B2(G210), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n541), .A2(new_n547), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(new_n545), .Z(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n863), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n868), .B2(new_n872), .ZN(G51));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n864), .B2(new_n865), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n854), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n717), .B(KEYINPUT57), .Z(new_n878));
  OAI22_X1  g692(.A1(new_n877), .A2(new_n878), .B1(new_n597), .B2(new_n596), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n867), .A2(new_n746), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n862), .B1(new_n879), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n867), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n882), .A2(KEYINPUT122), .A3(new_n462), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n863), .B1(new_n882), .B2(new_n462), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n882), .B2(new_n462), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G60));
  AND2_X1   g700(.A1(new_n618), .A2(new_n620), .ZN(new_n887));
  NAND2_X1  g701(.A1(G478), .A2(G902), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT59), .Z(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n862), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n850), .B2(new_n854), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(new_n887), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n892), .C1(new_n893), .C2(new_n887), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT60), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n866), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n642), .B2(new_n641), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n370), .B(new_n371), .C1(new_n866), .C2(new_n900), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n863), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n902), .A2(KEYINPUT61), .A3(new_n863), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(G66));
  INV_X1    g722(.A(new_n483), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n272), .B1(new_n909), .B2(new_n516), .ZN(new_n910));
  INV_X1    g724(.A(new_n845), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n272), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n869), .B1(G898), .B2(new_n272), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n912), .B(new_n913), .Z(G69));
  OAI21_X1  g728(.A(new_n295), .B1(new_n245), .B2(new_n244), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n453), .B1(KEYINPUT19), .B2(new_n340), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT124), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n915), .B(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n757), .A2(new_n763), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n815), .A2(new_n711), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n750), .A2(new_n699), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n736), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n919), .A2(new_n741), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n272), .B1(new_n923), .B2(new_n738), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n272), .A2(G900), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n918), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n920), .A2(new_n670), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT62), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n928), .A2(KEYINPUT62), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n806), .B(KEYINPUT125), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n663), .A2(new_n719), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(new_n323), .A3(new_n385), .A4(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n919), .A2(new_n929), .A3(new_n930), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n272), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n918), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n927), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n927), .B2(new_n936), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G72));
  XOR2_X1   g754(.A(new_n657), .B(KEYINPUT63), .Z(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n934), .B2(new_n911), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n264), .A2(new_n290), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n276), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n862), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n941), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n923), .A2(new_n738), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n845), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n276), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n279), .A2(new_n286), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n951), .B2(new_n316), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n838), .B2(new_n849), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(G57));
endmodule


