//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G110), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n196), .C1(new_n191), .C2(G128), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(new_n194), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n195), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT24), .B(G110), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT73), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(new_n206), .A3(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT16), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n210), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G146), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT66), .A2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT66), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G125), .B(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n207), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n212), .A2(new_n213), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT72), .A3(new_n214), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n201), .A2(new_n202), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G110), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT74), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT74), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G137), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n236), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n239), .B(KEYINPUT75), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n221), .A2(new_n231), .A3(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n188), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT76), .B(KEYINPUT25), .Z(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(KEYINPUT25), .A3(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n246), .B2(new_n248), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n189), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n189), .A2(G902), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n242), .A2(new_n243), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G472), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT66), .A2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT66), .A2(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(G143), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n260), .A2(new_n266), .A3(new_n261), .A4(new_n263), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n262), .A2(G146), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n217), .B2(G143), .ZN(new_n270));
  OR3_X1    g084(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n261), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n265), .A2(new_n267), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(G137), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(KEYINPUT68), .A2(G131), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(G134), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n280), .A3(G131), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n260), .A2(new_n263), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n199), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n258), .A2(new_n259), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n268), .B1(new_n292), .B2(new_n262), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n274), .A2(new_n283), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT2), .B(G113), .Z(new_n298));
  XNOR2_X1  g112(.A(G116), .B(G119), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n191), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n297), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n299), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n305), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n295), .A2(new_n296), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n265), .A2(new_n267), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n270), .A2(new_n273), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n283), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n294), .A2(new_n288), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n311), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n288), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n294), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n315), .ZN(new_n324));
  INV_X1    g138(.A(new_n311), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(G237), .A2(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G210), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT27), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G101), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n315), .A2(KEYINPUT30), .A3(new_n316), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n217), .B2(G143), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n270), .B1(new_n336), .B2(new_n199), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n337), .A2(new_n290), .B1(new_n288), .B2(new_n320), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n338), .A2(new_n322), .B1(new_n274), .B2(new_n283), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n325), .B(new_n334), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(new_n317), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n332), .B(new_n333), .C1(new_n343), .C2(new_n331), .ZN(new_n344));
  INV_X1    g158(.A(new_n295), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n312), .A2(new_n318), .B1(new_n325), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n331), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n333), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n257), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n317), .A3(new_n331), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n342), .A2(KEYINPUT31), .A3(new_n317), .A4(new_n331), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n319), .A2(new_n326), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n347), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n350), .B1(new_n359), .B2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n356), .B2(new_n358), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n256), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n237), .A2(G952), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(G237), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT21), .B(G898), .Z(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT91), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n188), .B(new_n237), .C1(G234), .C2(G237), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT7), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n237), .A2(G224), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT82), .Z(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n313), .A2(G125), .A3(new_n314), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n294), .A2(new_n210), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n374), .B(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(G113), .B1(new_n301), .B2(KEYINPUT5), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(KEYINPUT5), .B2(new_n299), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n306), .ZN(new_n385));
  OR2_X1    g199(.A1(KEYINPUT78), .A2(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT78), .A2(G104), .ZN(new_n387));
  AOI21_X1  g201(.A(G107), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(G104), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT79), .A3(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n390), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n397), .A3(new_n387), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NOR2_X1   g213(.A1(KEYINPUT3), .A2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT3), .A2(G107), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n385), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(G110), .B(G122), .Z(new_n406));
  XOR2_X1   g220(.A(new_n406), .B(KEYINPUT8), .Z(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n383), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT83), .B(G113), .C1(new_n301), .C2(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n412), .A2(new_n308), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n405), .B(new_n407), .C1(new_n413), .C2(new_n404), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n373), .B1(new_n380), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n378), .A2(new_n379), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT7), .A3(new_n376), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT84), .A3(new_n382), .A4(new_n414), .ZN(new_n419));
  INV_X1    g233(.A(new_n387), .ZN(new_n420));
  NOR2_X1   g234(.A1(KEYINPUT78), .A2(G104), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n420), .A2(new_n400), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n402), .B1(new_n397), .B2(new_n392), .ZN(new_n423));
  OAI21_X1  g237(.A(G101), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(G101), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n310), .A3(new_n307), .A4(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n406), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n395), .A2(new_n403), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n385), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n419), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n417), .A2(new_n376), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n378), .A2(new_n377), .A3(new_n379), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n406), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  AND4_X1   g255(.A1(new_n440), .A2(new_n437), .A3(new_n441), .A4(new_n406), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n429), .B1(new_n428), .B2(new_n431), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n443), .B2(new_n441), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n436), .B(new_n439), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n433), .A2(new_n445), .A3(new_n188), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n433), .A2(new_n445), .A3(new_n188), .A4(new_n447), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n370), .B(new_n372), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT9), .B(G234), .ZN(new_n452));
  OAI21_X1  g266(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n237), .A2(G227), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n283), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT10), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n404), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n260), .A2(new_n263), .A3(new_n289), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT1), .B1(new_n262), .B2(G146), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n260), .A2(new_n263), .B1(G128), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n403), .B(new_n395), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n460), .A2(new_n294), .B1(new_n464), .B2(new_n459), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n313), .A2(new_n425), .A3(new_n314), .A4(new_n427), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n459), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n430), .A2(KEYINPUT10), .A3(new_n294), .ZN(new_n469));
  AND4_X1   g283(.A1(new_n458), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n457), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n466), .A2(new_n469), .A3(new_n468), .A4(new_n458), .ZN(new_n472));
  INV_X1    g286(.A(new_n457), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n464), .B1(new_n430), .B2(new_n294), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n474), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT12), .B1(new_n474), .B2(new_n283), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n472), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(G469), .B(G902), .C1(new_n471), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G469), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n188), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(new_n283), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(KEYINPUT12), .A3(new_n283), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n473), .B1(new_n486), .B2(new_n472), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n467), .A2(new_n470), .A3(new_n457), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT80), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n475), .A2(new_n476), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n457), .B1(new_n490), .B2(new_n470), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n492));
  INV_X1    g306(.A(new_n467), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n472), .A3(new_n473), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n495), .A3(G469), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n454), .B1(new_n481), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  NOR2_X1   g312(.A1(G475), .A2(G902), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n392), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n327), .A2(G143), .A3(G214), .ZN(new_n502));
  AOI21_X1  g316(.A(G143), .B1(new_n327), .B2(G214), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n237), .A3(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n262), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n327), .A2(G143), .A3(G214), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(KEYINPUT86), .A3(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n284), .A3(new_n510), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n512), .A3(new_n516), .A4(new_n513), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n218), .B1(KEYINPUT88), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n218), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n214), .B1(new_n521), .B2(new_n292), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n209), .A2(new_n211), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G146), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n526), .A2(KEYINPUT85), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n219), .B1(new_n526), .B2(KEYINPUT85), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n511), .A2(KEYINPUT18), .A3(G131), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n509), .A2(new_n510), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n501), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n225), .A2(new_n227), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT86), .B1(new_n511), .B2(G131), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n505), .B(new_n284), .C1(new_n509), .C2(new_n510), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT17), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n506), .A2(new_n512), .A3(new_n540), .A4(new_n513), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n542), .A2(new_n534), .A3(new_n501), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n498), .B(new_n499), .C1(new_n535), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n535), .A2(new_n543), .ZN(new_n546));
  INV_X1    g360(.A(new_n499), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT20), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n534), .A3(new_n501), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n529), .A2(new_n533), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n522), .B1(KEYINPUT87), .B2(new_n514), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n517), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n549), .B1(new_n552), .B2(new_n501), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n498), .A4(new_n499), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n557));
  XNOR2_X1  g371(.A(G116), .B(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n390), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n262), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n199), .A2(G143), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n276), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n276), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n559), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n302), .A2(KEYINPUT14), .A3(G122), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G107), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT14), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(new_n558), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n557), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(G116), .B(G122), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G107), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n563), .B1(new_n572), .B2(new_n559), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT13), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n560), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n561), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n560), .A2(new_n574), .ZN(new_n577));
  OAI21_X1  g391(.A(G134), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(G107), .B(new_n566), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n560), .A2(new_n561), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G134), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n562), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n580), .A2(new_n583), .A3(KEYINPUT90), .A4(new_n559), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n570), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n452), .A2(new_n187), .A3(G953), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n580), .A2(new_n583), .A3(new_n559), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(new_n557), .B1(new_n573), .B2(new_n578), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n584), .A3(new_n586), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n592), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n501), .B1(new_n542), .B2(new_n534), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n188), .B1(new_n543), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G475), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n556), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n497), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n363), .A2(new_n451), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  AND3_X1   g418(.A1(new_n497), .A2(new_n253), .A3(new_n255), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n356), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n353), .A2(new_n354), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n355), .A2(new_n347), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n357), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n556), .A2(new_n600), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n585), .A2(new_n587), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n586), .B1(new_n590), .B2(new_n584), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n188), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT93), .A3(new_n593), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT93), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n592), .B2(G478), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT33), .B1(new_n616), .B2(new_n617), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n588), .A2(new_n591), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n593), .A2(G902), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n619), .A2(new_n621), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT94), .B1(new_n615), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n630), .B(new_n627), .C1(new_n556), .C2(new_n600), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n451), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n451), .B(KEYINPUT95), .C1(new_n629), .C2(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n614), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AOI21_X1  g454(.A(new_n372), .B1(new_n449), .B2(new_n450), .ZN(new_n641));
  INV_X1    g455(.A(new_n370), .ZN(new_n642));
  INV_X1    g456(.A(new_n544), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n498), .B1(new_n553), .B2(new_n499), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n596), .B(new_n600), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n451), .A2(KEYINPUT97), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n614), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  INV_X1    g469(.A(new_n254), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n221), .A2(new_n234), .A3(new_n231), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n234), .B1(new_n221), .B2(new_n231), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n656), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n657), .A2(new_n658), .A3(new_n240), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n248), .B1(new_n664), .B2(new_n244), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT77), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n250), .A3(new_n249), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n663), .B1(new_n667), .B2(new_n189), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n655), .B1(new_n611), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n663), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n253), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(KEYINPUT98), .A3(new_n610), .A4(new_n606), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n602), .A3(new_n672), .A4(new_n451), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n449), .A2(new_n450), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n371), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n668), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n365), .B1(new_n369), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n645), .B2(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n548), .A2(new_n544), .B1(G475), .B2(new_n599), .ZN(new_n683));
  INV_X1    g497(.A(new_n681), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(KEYINPUT99), .A3(new_n596), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n609), .A2(KEYINPUT32), .A3(new_n357), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n344), .A2(new_n349), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G472), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n362), .A3(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n678), .A2(new_n686), .A3(new_n690), .A4(new_n497), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n676), .B(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n597), .B1(new_n556), .B2(new_n600), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n371), .A2(new_n695), .A3(new_n668), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n345), .A2(new_n325), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n331), .B1(new_n698), .B2(new_n317), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n343), .B2(new_n331), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n687), .A2(new_n362), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n687), .A2(new_n362), .A3(KEYINPUT101), .A4(new_n701), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n681), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n497), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND3_X1  g523(.A1(new_n697), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NAND3_X1  g525(.A1(new_n615), .A2(new_n628), .A3(new_n684), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n678), .A2(new_n690), .A3(new_n497), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  INV_X1    g529(.A(new_n256), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n471), .A2(new_n477), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n479), .B1(new_n717), .B2(new_n188), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n478), .A3(new_n454), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n716), .A2(new_n690), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n634), .B2(new_n635), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT41), .B(G113), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT102), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  AOI21_X1  g538(.A(new_n720), .B1(new_n650), .B2(new_n649), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n302), .ZN(G18));
  NAND2_X1  g540(.A1(new_n717), .A2(new_n188), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n479), .A3(new_n188), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n642), .A3(new_n453), .A4(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n596), .A3(new_n615), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n690), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n671), .A2(new_n641), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT103), .B(G119), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G21));
  INV_X1    g550(.A(new_n346), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n347), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n358), .B1(new_n607), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n609), .A2(new_n188), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(G472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n716), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n641), .A2(new_n642), .A3(new_n696), .A4(new_n719), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(G122), .Z(G24));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  AOI21_X1  g561(.A(G902), .B1(new_n607), .B2(new_n608), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n353), .A2(new_n354), .B1(new_n347), .B2(new_n737), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n748), .A2(new_n257), .B1(new_n358), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n750), .B2(new_n668), .ZN(new_n751));
  INV_X1    g565(.A(new_n739), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n671), .A2(KEYINPUT104), .A3(new_n606), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n627), .B1(new_n556), .B2(new_n600), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n641), .A2(new_n755), .A3(new_n684), .A4(new_n719), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n746), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g572(.A(KEYINPUT105), .B(new_n756), .C1(new_n751), .C2(new_n753), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n210), .ZN(G27));
  INV_X1    g575(.A(new_n480), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n491), .A2(new_n494), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n729), .B(new_n762), .C1(new_n479), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n453), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n449), .A2(new_n371), .A3(new_n450), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n712), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT106), .B(new_n361), .C1(new_n356), .C2(new_n358), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n362), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n360), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(KEYINPUT107), .A3(new_n716), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT107), .B1(new_n772), .B2(new_n716), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n765), .A2(new_n766), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n363), .A2(new_n713), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT108), .B(G131), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G33));
  NAND3_X1  g596(.A1(new_n363), .A2(new_n686), .A3(new_n776), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n763), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n489), .A2(new_n495), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n479), .B1(new_n787), .B2(new_n785), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n788), .B2(KEYINPUT109), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(KEYINPUT109), .B2(new_n788), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT110), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT46), .B1(new_n790), .B2(new_n762), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n478), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n454), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n707), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n628), .A2(new_n556), .A3(new_n600), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT43), .Z(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n611), .A3(new_n671), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n799), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n766), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n799), .B2(new_n800), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT111), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT112), .B(G137), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G39));
  NOR4_X1   g622(.A1(new_n716), .A2(new_n690), .A3(new_n712), .A4(new_n766), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n811), .B(new_n454), .C1(new_n792), .C2(new_n794), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NOR2_X1   g628(.A1(new_n718), .A2(new_n478), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n372), .B(new_n454), .C1(new_n816), .C2(KEYINPUT49), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(KEYINPUT49), .B2(new_n816), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n695), .A3(new_n797), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n706), .A2(new_n256), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n716), .A2(new_n798), .A3(new_n365), .A4(new_n741), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n719), .A2(new_n372), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT117), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n694), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n802), .A2(new_n365), .A3(new_n719), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n828), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n829), .A2(new_n615), .A3(new_n628), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n798), .A2(new_n828), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n754), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n816), .A2(new_n453), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n810), .A2(new_n812), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n822), .A2(new_n802), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n719), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n677), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n364), .B1(new_n822), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n629), .A2(new_n631), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n829), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n773), .A2(new_n774), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT118), .A3(KEYINPUT48), .A4(new_n832), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n832), .ZN(new_n849));
  XOR2_X1   g663(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n850));
  AOI211_X1 g664(.A(new_n845), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n810), .ZN(new_n852));
  INV_X1    g666(.A(new_n812), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n837), .B(KEYINPUT116), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n839), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n834), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n840), .B(new_n851), .C1(new_n857), .C2(KEYINPUT51), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n704), .A2(new_n705), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n764), .A2(new_n453), .A3(new_n684), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n641), .A3(new_n668), .A4(new_n696), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n691), .B(new_n714), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n760), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT104), .B1(new_n741), .B2(new_n671), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n750), .A2(new_n747), .A3(new_n668), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n757), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT105), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n754), .A2(new_n746), .A3(new_n757), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n691), .A2(new_n714), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n862), .B1(new_n704), .B2(new_n705), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n754), .A2(new_n767), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n690), .A2(new_n497), .A3(new_n671), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n449), .A2(new_n450), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n618), .A2(new_n594), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n592), .A2(new_n595), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n681), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n600), .C1(new_n643), .C2(new_n644), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n878), .A2(new_n883), .A3(new_n884), .A4(new_n371), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT113), .B1(new_n766), .B2(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n877), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n876), .A2(new_n783), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n601), .B1(new_n615), .B2(new_n627), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n605), .A2(new_n451), .A3(new_n890), .A4(new_n612), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n673), .A3(new_n603), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n732), .A2(new_n733), .B1(new_n742), .B2(new_n743), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n721), .A2(new_n725), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n893), .A2(new_n895), .A3(new_n780), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n875), .A2(new_n896), .A3(KEYINPUT53), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n875), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n760), .A2(new_n859), .A3(new_n863), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT52), .B1(new_n870), .B2(new_n873), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n893), .A2(new_n895), .A3(new_n780), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n875), .A2(new_n896), .A3(KEYINPUT53), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n905), .A2(KEYINPUT115), .A3(new_n906), .A4(new_n907), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n858), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n821), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n237), .A2(G952), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n436), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n905), .A2(new_n906), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  INV_X1    g734(.A(G210), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(KEYINPUT119), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n918), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n918), .A2(KEYINPUT120), .ZN(new_n927));
  OAI221_X1 g741(.A(new_n924), .B1(KEYINPUT119), .B2(new_n927), .C1(new_n920), .C2(new_n921), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n915), .B1(new_n926), .B2(new_n928), .ZN(G51));
  XNOR2_X1  g743(.A(new_n919), .B(new_n907), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n480), .B(KEYINPUT57), .Z(new_n931));
  OAI21_X1  g745(.A(new_n717), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n920), .A2(new_n790), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n915), .B1(new_n932), .B2(new_n933), .ZN(G54));
  NAND4_X1  g748(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n546), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n546), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n915), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n910), .A2(new_n911), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n625), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT121), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  INV_X1    g759(.A(new_n915), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n625), .A2(new_n941), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n930), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(new_n661), .A2(new_n662), .ZN(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND3_X1  g766(.A1(new_n919), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n950), .A4(new_n952), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n946), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n897), .B2(new_n898), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n242), .A2(new_n243), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G66));
  INV_X1    g777(.A(G224), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n368), .B2(new_n964), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n892), .A2(new_n721), .A3(new_n725), .A4(new_n894), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n916), .B1(G898), .B2(new_n237), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n967), .B(new_n969), .ZN(G69));
  AOI22_X1  g784(.A1(new_n324), .A2(new_n340), .B1(new_n295), .B2(KEYINPUT30), .ZN(new_n971));
  INV_X1    g785(.A(new_n521), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(G900), .B2(G953), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n641), .A2(new_n696), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n796), .A2(new_n978), .A3(new_n846), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n760), .A2(new_n871), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n980), .A2(new_n780), .A3(new_n783), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n806), .A2(new_n979), .A3(new_n813), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n976), .B1(new_n982), .B2(new_n237), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n710), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  INV_X1    g799(.A(new_n708), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n363), .A2(new_n986), .A3(new_n802), .A4(new_n890), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n796), .B2(new_n805), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n989), .A3(new_n813), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n973), .B1(new_n990), .B2(new_n237), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n983), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n237), .B1(G227), .B2(G900), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n994), .C1(new_n983), .C2(new_n991), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  XNOR2_X1  g812(.A(new_n343), .B(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n347), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n982), .A2(new_n966), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n985), .A2(new_n989), .A3(new_n813), .A4(new_n966), .ZN(new_n1005));
  AOI211_X1 g819(.A(new_n347), .B(new_n999), .C1(new_n1005), .C2(new_n1003), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n343), .B(new_n331), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n905), .B2(new_n906), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1004), .A2(new_n1006), .A3(new_n915), .A4(new_n1010), .ZN(G57));
endmodule


