//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n460), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n469), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n468), .B1(new_n477), .B2(G2105), .ZN(G160));
  INV_X1    g053(.A(new_n466), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT68), .Z(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n463), .B1(new_n471), .B2(new_n473), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT69), .Z(new_n490));
  AND3_X1   g065(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n469), .A2(new_n474), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n501), .A3(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT5), .B1(new_n511), .B2(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  INV_X1    g098(.A(new_n517), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n510), .A2(new_n514), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n529), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n525), .A2(new_n527), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(G52), .A2(new_n524), .B1(new_n526), .B2(G90), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n521), .B2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G43), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n524), .A2(new_n538), .B1(new_n526), .B2(G81), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n521), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n524), .A2(G53), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n515), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n551), .B(new_n554), .C1(new_n521), .C2(new_n555), .ZN(G299));
  INV_X1    g131(.A(G166), .ZN(G303));
  NAND2_X1  g132(.A1(new_n526), .A2(new_n552), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G87), .A3(new_n559), .ZN(new_n560));
  OR3_X1    g135(.A1(new_n512), .A2(new_n513), .A3(G74), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n524), .A2(G49), .B1(G651), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(G288));
  NOR2_X1   g138(.A1(new_n512), .A2(new_n513), .ZN(new_n564));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT74), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G73), .ZN(new_n567));
  INV_X1    g142(.A(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g144(.A1(new_n564), .A2(KEYINPUT74), .A3(new_n565), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n553), .A2(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  AOI22_X1  g149(.A1(G47), .A2(new_n524), .B1(new_n526), .B2(G85), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n521), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n553), .A2(G92), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT75), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n585));
  INV_X1    g160(.A(G54), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n586), .B1(new_n517), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT77), .B1(new_n589), .B2(new_n568), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n589), .A2(new_n568), .A3(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n564), .C2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n585), .A2(new_n588), .B1(G651), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n583), .A2(new_n584), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n579), .B1(new_n595), .B2(G868), .ZN(G321));
  XNOR2_X1  g171(.A(G321), .B(KEYINPUT78), .ZN(G284));
  MUX2_X1   g172(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n595), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g180(.A1(new_n469), .A2(new_n474), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n461), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n488), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n463), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G135), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n614), .B1(new_n615), .B2(new_n616), .C1(new_n482), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n631), .ZN(G401));
  XOR2_X1   g212(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  INV_X1    g220(.A(new_n638), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  AOI211_X1 g234(.A(new_n657), .B(new_n659), .C1(new_n652), .C2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  XOR2_X1   g237(.A(G1991), .B(G1996), .Z(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT82), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(G229));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G20), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT23), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(G299), .B2(G16), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G1956), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n543), .A2(new_n670), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(G19), .ZN(new_n676));
  INV_X1    g251(.A(G1341), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n618), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT92), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G11), .ZN(new_n682));
  AND2_X1   g257(.A1(KEYINPUT30), .A2(G28), .ZN(new_n683));
  NOR2_X1   g258(.A1(KEYINPUT30), .A2(G28), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G1961), .ZN(new_n687));
  NOR2_X1   g262(.A1(G171), .A2(new_n670), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G5), .B2(new_n670), .ZN(new_n689));
  AOI211_X1 g264(.A(new_n678), .B(new_n686), .C1(new_n687), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n679), .A2(G32), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n483), .A2(G141), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n461), .A2(G105), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT26), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n693), .B(new_n695), .C1(G129), .C2(new_n488), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n691), .B1(new_n698), .B2(new_n679), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT27), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n679), .A2(G26), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n488), .A2(G128), .ZN(new_n704));
  NOR2_X1   g279(.A1(G104), .A2(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT88), .Z(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n707));
  INV_X1    g282(.A(G140), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n704), .B1(new_n706), .B2(new_n707), .C1(new_n482), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(G29), .ZN(new_n710));
  INV_X1    g285(.A(G2067), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  NAND2_X1  g289(.A1(G168), .A2(G16), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(KEYINPUT90), .C1(G16), .C2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(KEYINPUT90), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT91), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n690), .B(new_n713), .C1(new_n714), .C2(new_n718), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n674), .B(new_n719), .C1(new_n714), .C2(new_n718), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n689), .A2(new_n687), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n679), .B1(new_n723), .B2(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G160), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2084), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n679), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n679), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2078), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n679), .A2(G33), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n606), .A2(G127), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n463), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT89), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI211_X1 g313(.A(new_n735), .B(new_n738), .C1(G139), .C2(new_n483), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n679), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2072), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n731), .B(new_n741), .C1(new_n677), .C2(new_n676), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G35), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G162), .B2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n728), .B(new_n742), .C1(new_n746), .C2(G2090), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G2090), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n670), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n595), .B2(new_n670), .ZN(new_n750));
  INV_X1    g325(.A(G1348), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n720), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G6), .B(G305), .S(G16), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G23), .ZN(new_n757));
  NAND2_X1  g332(.A1(G288), .A2(KEYINPUT85), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n560), .A2(new_n759), .A3(new_n562), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n757), .B1(new_n761), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT33), .B(G1976), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n670), .A2(G22), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G166), .B2(new_n670), .ZN(new_n766));
  INV_X1    g341(.A(G1971), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n756), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT34), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT86), .Z(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(KEYINPUT34), .ZN(new_n772));
  NOR2_X1   g347(.A1(G25), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n483), .A2(G131), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n775));
  INV_X1    g350(.A(G107), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G2105), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G119), .B2(new_n488), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n773), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT35), .B(G1991), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT83), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n781), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G290), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G16), .B2(G24), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT84), .B(G1986), .Z(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n772), .A2(new_n784), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n771), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n771), .A2(KEYINPUT36), .A3(new_n792), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n753), .A2(new_n795), .A3(new_n796), .ZN(G311));
  INV_X1    g372(.A(G311), .ZN(G150));
  NAND2_X1  g373(.A1(new_n595), .A2(G559), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT38), .ZN(new_n800));
  AOI22_X1  g375(.A1(G55), .A2(new_n524), .B1(new_n526), .B2(G93), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n521), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n543), .B(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n800), .B(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT39), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(KEYINPUT39), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n806), .A2(new_n807), .A3(G860), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n803), .A2(G860), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT37), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n810), .ZN(G145));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n739), .B2(KEYINPUT96), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n812), .B2(new_n739), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n697), .B(new_n709), .Z(new_n815));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n498), .A2(new_n816), .A3(new_n502), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n498), .B2(new_n502), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n497), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(new_n814), .B(new_n813), .S(new_n820), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n779), .B(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n488), .A2(G130), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G118), .B2(new_n463), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n483), .B2(G142), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n609), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n821), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n618), .B(G160), .Z(new_n833));
  XNOR2_X1  g408(.A(G162), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n832), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT100), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g413(.A1(new_n803), .A2(G868), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n595), .A2(G299), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n595), .A2(G299), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n595), .A2(KEYINPUT101), .A3(G299), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n602), .B(new_n804), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(KEYINPUT41), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n840), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n761), .B(new_n785), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G305), .B(G303), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT42), .Z(new_n860));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n847), .B1(new_n851), .B2(new_n846), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n861), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  AOI21_X1  g439(.A(new_n839), .B1(new_n864), .B2(G868), .ZN(G295));
  AOI21_X1  g440(.A(new_n839), .B1(new_n864), .B2(G868), .ZN(G331));
  XNOR2_X1  g441(.A(new_n804), .B(G301), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G286), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n845), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n851), .B2(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n859), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  INV_X1    g449(.A(new_n859), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n868), .B1(new_n848), .B2(new_n850), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n870), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT44), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n868), .A2(new_n849), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n840), .A2(new_n842), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n859), .B(new_n882), .C1(new_n845), .C2(new_n880), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n874), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n877), .A2(new_n886), .A3(new_n874), .A4(new_n883), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(KEYINPUT43), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n879), .A2(new_n888), .A3(KEYINPUT105), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT105), .B1(new_n879), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n872), .A2(new_n874), .A3(new_n877), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(KEYINPUT43), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n889), .A2(new_n890), .B1(KEYINPUT44), .B2(new_n893), .ZN(G397));
  NAND2_X1  g469(.A1(new_n503), .A2(KEYINPUT95), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n498), .A2(new_n816), .A3(new_n502), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G1384), .B1(new_n897), .B2(new_n497), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT50), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G1384), .B1(new_n497), .B2(new_n504), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n477), .A2(G2105), .ZN(new_n904));
  INV_X1    g479(.A(new_n468), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G40), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(G2084), .ZN(new_n909));
  INV_X1    g484(.A(new_n898), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n901), .A2(KEYINPUT45), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n714), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(G8), .B1(new_n916), .B2(G286), .ZN(new_n917));
  AOI21_X1  g492(.A(G168), .B1(new_n909), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT51), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(KEYINPUT51), .B2(new_n917), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n922));
  OAI211_X1 g497(.A(G160), .B(G40), .C1(new_n901), .C2(KEYINPUT45), .ZN(new_n923));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n819), .A2(KEYINPUT45), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT109), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n819), .A2(new_n927), .A3(KEYINPUT45), .A4(new_n924), .ZN(new_n928));
  AOI211_X1 g503(.A(new_n922), .B(new_n923), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(new_n923), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT110), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n921), .B1(new_n933), .B2(G2078), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n908), .A2(new_n687), .ZN(new_n935));
  XOR2_X1   g510(.A(G301), .B(KEYINPUT54), .Z(new_n936));
  NAND2_X1  g511(.A1(new_n912), .A2(new_n907), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(new_n938), .A3(G2078), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n930), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n940), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n939), .A2(new_n913), .B1(new_n687), .B2(new_n908), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT124), .Z(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n934), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n920), .B(new_n941), .C1(new_n944), .C2(new_n936), .ZN(new_n945));
  XOR2_X1   g520(.A(G299), .B(KEYINPUT57), .Z(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n927), .B1(new_n898), .B2(KEYINPUT45), .ZN(new_n948));
  INV_X1    g523(.A(new_n928), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n931), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(G2072), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1956), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n907), .B1(KEYINPUT50), .B2(new_n902), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n898), .A2(new_n899), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n959), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n960), .A2(KEYINPUT121), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(KEYINPUT120), .A2(KEYINPUT61), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n960), .B2(new_n962), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n946), .A2(new_n961), .A3(KEYINPUT121), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT61), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n910), .A2(new_n906), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT58), .B(G1341), .Z(new_n972));
  AOI22_X1  g547(.A1(new_n951), .A2(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(new_n542), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n908), .A2(new_n751), .B1(new_n970), .B2(new_n711), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n595), .A2(new_n977), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(KEYINPUT123), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n583), .A2(new_n584), .A3(new_n594), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(KEYINPUT60), .A3(new_n976), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT122), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT122), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(KEYINPUT123), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n979), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT120), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n968), .B(new_n987), .C1(new_n988), .C2(new_n965), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n960), .A2(new_n980), .A3(new_n976), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n962), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n945), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n572), .A2(new_n993), .A3(new_n573), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n526), .A2(G86), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n572), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT49), .B(new_n994), .C1(new_n996), .C2(new_n993), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n572), .A2(new_n993), .A3(new_n573), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n572), .B2(new_n995), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n970), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n758), .A2(G1976), .A3(new_n760), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n758), .A2(new_n1007), .A3(G1976), .A4(new_n760), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1006), .A2(new_n1003), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1004), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n950), .A2(new_n922), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n930), .A2(KEYINPUT110), .A3(new_n931), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n767), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n908), .A2(G2090), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  OAI22_X1  g595(.A1(G166), .A2(new_n1002), .B1(KEYINPUT111), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1019), .A2(KEYINPUT112), .A3(G8), .A4(new_n1023), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1023), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n956), .A2(G2090), .A3(new_n957), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n933), .B2(new_n767), .ZN(new_n1031));
  OAI211_X1 g606(.A(KEYINPUT114), .B(new_n1029), .C1(new_n1031), .C2(new_n1002), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1002), .B1(new_n1017), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(new_n1023), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n992), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1004), .A2(new_n1011), .A3(new_n560), .A4(new_n562), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1003), .B1(new_n1042), .B2(new_n999), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n1014), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n916), .A2(G8), .A3(G168), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(KEYINPUT63), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1019), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(new_n1028), .C1(new_n1023), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1014), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1044), .A2(new_n1037), .A3(new_n1054), .A4(new_n1048), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT116), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1028), .A2(new_n1058), .A3(new_n1037), .A4(new_n1048), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1056), .A2(KEYINPUT117), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1063));
  AOI211_X1 g638(.A(KEYINPUT118), .B(new_n1045), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1055), .A2(KEYINPUT116), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n1057), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n1063), .A3(new_n1052), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1045), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1040), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT127), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT127), .B(new_n1040), .C1(new_n1064), .C2(new_n1071), .ZN(new_n1075));
  AOI211_X1 g650(.A(G301), .B(new_n944), .C1(KEYINPUT62), .C2(new_n920), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n1039), .C1(KEYINPUT62), .C2(new_n920), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n779), .B(new_n782), .ZN(new_n1079));
  XOR2_X1   g654(.A(new_n1079), .B(KEYINPUT108), .Z(new_n1080));
  XNOR2_X1  g655(.A(new_n709), .B(new_n711), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n698), .A2(G1996), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n697), .A2(new_n969), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G290), .A2(G1986), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT107), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(G1986), .B2(G290), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT106), .B1(new_n912), .B2(new_n906), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1078), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(KEYINPUT48), .A3(new_n1087), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT48), .B1(new_n1093), .B2(new_n1087), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT46), .B1(new_n1093), .B2(new_n969), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n698), .B2(new_n1081), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT46), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1092), .A2(new_n1102), .A3(G1996), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT47), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n780), .A2(new_n782), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1084), .A2(new_n1106), .B1(G2067), .B2(new_n709), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1099), .B(new_n1105), .C1(new_n1093), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g684(.A(G319), .ZN(new_n1111));
  NOR3_X1   g685(.A1(G401), .A2(new_n1111), .A3(G227), .ZN(new_n1112));
  NAND4_X1  g686(.A1(new_n837), .A2(new_n668), .A3(new_n667), .A4(new_n1112), .ZN(new_n1113));
  NOR2_X1   g687(.A1(new_n1113), .A2(new_n893), .ZN(G308));
  INV_X1    g688(.A(G308), .ZN(G225));
endmodule


