//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n208), .B1(new_n209), .B2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT1), .B1(new_n211), .B2(G127gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(G134gat), .ZN(new_n213));
  XOR2_X1   g012(.A(KEYINPUT69), .B(G134gat), .Z(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n209), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  INV_X1    g015(.A(new_n208), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n207), .A2(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n210), .A2(new_n212), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G155gat), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G148gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT74), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT74), .B1(new_n228), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(G162gat), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT75), .B1(new_n236), .B2(KEYINPUT2), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n230), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT75), .B1(new_n223), .B2(new_n225), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n239), .B(new_n240), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n221), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n226), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n248), .A2(new_n249), .A3(new_n222), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n239), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n229), .A2(G148gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n227), .A2(G141gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n242), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT74), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(KEYINPUT77), .A3(new_n243), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n220), .B1(new_n245), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n243), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n220), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n204), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n245), .B2(new_n258), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n238), .B2(new_n244), .ZN(new_n269));
  INV_X1    g068(.A(new_n220), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n265), .B(new_n266), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n262), .A2(new_n203), .ZN(new_n273));
  OAI211_X1 g072(.A(KEYINPUT5), .B(new_n263), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n268), .A2(new_n271), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(new_n265), .A3(new_n266), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G57gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n274), .A2(new_n277), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G8gat), .B(G36gat), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(G64gat), .ZN(new_n289));
  INV_X1    g088(.A(G92gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT68), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  INV_X1    g099(.A(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n299), .B1(new_n304), .B2(KEYINPUT68), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n296), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  INV_X1    g107(.A(G183gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT27), .B1(new_n309), .B2(KEYINPUT66), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(G190gat), .ZN(new_n314));
  AND4_X1   g113(.A1(new_n308), .A2(new_n310), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n308), .B1(new_n316), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT67), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n312), .A2(new_n309), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n314), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT28), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n310), .A2(new_n313), .A3(new_n308), .A4(new_n314), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n295), .A2(KEYINPUT64), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT64), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT65), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT24), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n327), .A2(new_n329), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n295), .A2(new_n330), .ZN(new_n335));
  NOR2_X1   g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n297), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n338), .A2(KEYINPUT25), .A3(new_n303), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n303), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n335), .A2(new_n346), .A3(new_n336), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AOI211_X1 g148(.A(KEYINPUT29), .B(new_n294), .C1(new_n326), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(G211gat), .ZN(new_n352));
  INV_X1    g151(.A(G218gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n351), .B(new_n354), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n351), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n351), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n355), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n326), .A2(new_n294), .A3(new_n349), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n350), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n326), .A2(new_n349), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n293), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n326), .A2(new_n294), .A3(new_n349), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n292), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT37), .B1(new_n366), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n364), .B1(new_n350), .B2(new_n365), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT37), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n367), .A3(new_n371), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n292), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT38), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n282), .B1(new_n274), .B2(new_n277), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT6), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n366), .A2(new_n372), .A3(KEYINPUT37), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n291), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT38), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n287), .A2(new_n382), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n390), .B(G22gat), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  INV_X1    g192(.A(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n267), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n238), .A2(new_n244), .A3(new_n221), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT77), .B1(new_n257), .B2(new_n243), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n257), .B2(new_n243), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n364), .B1(new_n401), .B2(KEYINPUT29), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n367), .B1(new_n269), .B2(new_n369), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n367), .B2(new_n369), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n396), .B1(new_n405), .B2(new_n260), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n403), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n245), .B2(new_n258), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n395), .B1(new_n411), .B2(new_n404), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n402), .B(new_n396), .C1(new_n260), .C2(new_n405), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n392), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n408), .B1(new_n403), .B2(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n413), .A3(new_n410), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n391), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n376), .A2(new_n291), .A3(new_n378), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n292), .C1(new_n366), .C2(new_n372), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT40), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n272), .A2(new_n204), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n259), .A2(new_n204), .A3(new_n262), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n426), .A2(KEYINPUT39), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT39), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n272), .A2(new_n429), .A3(new_n204), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n282), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n425), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(KEYINPUT39), .A3(new_n427), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n433), .A2(KEYINPUT40), .A3(new_n282), .A4(new_n430), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n424), .A2(new_n284), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n389), .A2(new_n419), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n368), .A2(new_n270), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n326), .A2(new_n220), .A3(new_n349), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT34), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n326), .A2(new_n220), .A3(new_n349), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n220), .B1(new_n326), .B2(new_n349), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n447), .B2(new_n441), .ZN(new_n448));
  NOR4_X1   g247(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT34), .A4(new_n442), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT72), .B(G15gat), .ZN(new_n455));
  INV_X1    g254(.A(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G71gat), .B(G99gat), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(new_n444), .A3(new_n441), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(KEYINPUT32), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n441), .A3(new_n439), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT34), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n450), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n450), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT36), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n284), .A2(KEYINPUT78), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n286), .A2(new_n285), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n383), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n424), .B1(new_n477), .B2(new_n384), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n436), .B(new_n472), .C1(new_n478), .C2(new_n419), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n460), .A3(new_n465), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n459), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n462), .A2(new_n461), .A3(new_n464), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n462), .B1(new_n464), .B2(new_n461), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND4_X1   g283(.A1(KEYINPUT35), .A2(new_n419), .A3(new_n480), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n286), .A2(new_n285), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n384), .B1(new_n486), .B2(new_n383), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n421), .A2(new_n423), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n468), .A3(new_n488), .A4(new_n419), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n478), .A2(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n202), .B1(new_n479), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n479), .A2(new_n202), .A3(new_n491), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT16), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(G1gat), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(G1gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(KEYINPUT83), .ZN(new_n501));
  NAND2_X1  g300(.A1(KEYINPUT84), .A2(G8gat), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n499), .A2(KEYINPUT84), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n502), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n498), .B1(KEYINPUT83), .B2(new_n504), .C1(G1gat), .C2(new_n496), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G8gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT14), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT80), .B(KEYINPUT15), .Z(new_n510));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n511));
  INV_X1    g310(.A(G50gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G43gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n456), .A2(KEYINPUT81), .A3(G50gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n514), .C1(new_n456), .C2(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n509), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT15), .B1(new_n456), .B2(G50gat), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n456), .B2(G50gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT82), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n518), .B1(new_n509), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT86), .B1(new_n507), .B2(new_n525), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT85), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT13), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n529), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n525), .B(KEYINPUT17), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n503), .A2(new_n506), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n526), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n531), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n535), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT11), .B(G169gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(G113gat), .B(G141gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n535), .A2(new_n542), .A3(new_n550), .A4(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT87), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n495), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OR3_X1    g357(.A1(new_n557), .A2(KEYINPUT88), .A3(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n507), .B1(KEYINPUT21), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n352), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(KEYINPUT21), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G127gat), .B(G155gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT20), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n566), .B(new_n568), .Z(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT19), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT89), .B(G183gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT7), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n575), .B(KEYINPUT91), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT8), .ZN(new_n582));
  NOR2_X1   g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(KEYINPUT92), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(new_n290), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n578), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT92), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n581), .A3(new_n587), .A4(new_n591), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n537), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  AND2_X1   g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n596), .A2(new_n525), .B1(KEYINPUT41), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G190gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n599), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n597), .A2(KEYINPUT41), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT90), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G218gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n596), .A2(new_n562), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n559), .B(new_n560), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n593), .A3(new_n594), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n301), .ZN(new_n616));
  INV_X1    g415(.A(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n608), .A2(new_n620), .A3(new_n610), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n562), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(KEYINPUT93), .A3(new_n622), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n614), .B(new_n619), .C1(new_n627), .C2(new_n613), .ZN(new_n628));
  INV_X1    g427(.A(new_n614), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n612), .B(KEYINPUT94), .Z(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n621), .B2(new_n622), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n618), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n574), .A2(new_n607), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n556), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n477), .A2(new_n384), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g441(.A1(new_n637), .A2(new_n488), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  AOI21_X1  g443(.A(KEYINPUT95), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT42), .ZN(new_n646));
  OAI21_X1  g445(.A(G8gat), .B1(new_n637), .B2(new_n488), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT96), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n638), .B2(new_n468), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT97), .ZN(new_n651));
  INV_X1    g450(.A(new_n472), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n638), .B2(new_n653), .ZN(G1326gat));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n419), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT43), .B(G22gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  INV_X1    g456(.A(new_n574), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n634), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n495), .A2(new_n555), .A3(new_n659), .A4(new_n607), .ZN(new_n660));
  INV_X1    g459(.A(G29gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n640), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT45), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n554), .A3(new_n634), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n493), .A2(KEYINPUT44), .A3(new_n494), .A4(new_n606), .ZN(new_n666));
  INV_X1    g465(.A(new_n384), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n383), .A2(new_n475), .ZN(new_n668));
  AOI211_X1 g467(.A(KEYINPUT78), .B(new_n282), .C1(new_n274), .C2(new_n277), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n668), .A2(new_n669), .A3(new_n486), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n485), .B(new_n488), .C1(new_n667), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n489), .A2(new_n490), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT99), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n675), .A2(new_n676), .B1(new_n677), .B2(new_n479), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n639), .A2(new_n488), .ZN(new_n679));
  INV_X1    g478(.A(new_n419), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n681), .A2(KEYINPUT98), .A3(new_n472), .A4(new_n436), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n607), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n665), .B(new_n666), .C1(new_n683), .C2(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n479), .A2(new_n677), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n491), .A2(KEYINPUT99), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT99), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n682), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n689), .B2(new_n606), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n665), .A4(new_n666), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n639), .B1(new_n685), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n663), .B1(new_n694), .B2(new_n661), .ZN(G1328gat));
  INV_X1    g494(.A(G36gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n660), .A2(new_n696), .A3(new_n424), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n685), .A2(new_n693), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n696), .B1(new_n699), .B2(new_n424), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n698), .B2(new_n700), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1329gat));
  OAI21_X1  g503(.A(G43gat), .B1(new_n684), .B2(new_n472), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n660), .A2(new_n456), .A3(new_n468), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n706), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n699), .A2(new_n652), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(G43gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n710), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n419), .B1(new_n685), .B2(new_n693), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n512), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n479), .A2(new_n202), .A3(new_n491), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n492), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n689), .A2(new_n606), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n692), .B1(new_n720), .B2(new_n665), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n690), .A2(new_n717), .A3(KEYINPUT100), .A4(new_n664), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n680), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n660), .A2(new_n512), .A3(new_n680), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n684), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(KEYINPUT103), .A3(new_n680), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G50gat), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT103), .B1(new_n729), .B2(new_n680), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT48), .B(new_n725), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n733), .ZN(G1331gat));
  NAND3_X1  g533(.A1(new_n574), .A2(new_n607), .A3(new_n633), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n554), .B(new_n735), .C1(new_n678), .C2(new_n682), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n640), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g537(.A(new_n488), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1333gat));
  AOI21_X1  g543(.A(G71gat), .B1(new_n736), .B2(new_n468), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n736), .A2(G71gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n652), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g547(.A1(new_n736), .A2(new_n680), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(new_n554), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n658), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n720), .A2(new_n633), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n639), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n718), .A2(new_n752), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(KEYINPUT106), .A3(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n639), .A2(G85gat), .A3(new_n634), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT107), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(G1336gat));
  OR2_X1    g564(.A1(new_n754), .A2(new_n488), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(new_n766), .B2(G92gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n633), .A2(new_n290), .A3(new_n424), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n758), .A2(new_n768), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(G92gat), .B2(new_n766), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n754), .B2(new_n472), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n760), .A2(new_n468), .A3(new_n761), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n634), .A2(G99gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(G1338gat));
  NOR3_X1   g576(.A1(new_n634), .A2(G106gat), .A3(new_n419), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT108), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n761), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n720), .A2(new_n680), .A3(new_n633), .A4(new_n753), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(KEYINPUT111), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n782), .B2(KEYINPUT111), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n780), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(G106gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n779), .B(KEYINPUT109), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n758), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT110), .B1(new_n789), .B2(KEYINPUT53), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n789), .A2(KEYINPUT110), .A3(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  NOR2_X1   g591(.A1(new_n635), .A2(new_n554), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n795));
  AOI21_X1  g594(.A(new_n619), .B1(new_n631), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n613), .B1(new_n625), .B2(new_n626), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n621), .A2(new_n622), .A3(new_n630), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT54), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT55), .B(new_n796), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n628), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n628), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n802), .A2(new_n554), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n540), .A2(KEYINPUT114), .A3(new_n541), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n543), .B2(new_n531), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n534), .B1(new_n529), .B2(new_n530), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n549), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n553), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n633), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n808), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n607), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  INV_X1    g621(.A(new_n807), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(KEYINPUT113), .B2(new_n801), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n606), .A3(new_n815), .A4(new_n804), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n658), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n822), .B1(new_n821), .B2(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n794), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n468), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n680), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n424), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n640), .A3(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT117), .Z(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n207), .A3(new_n554), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n834), .B2(new_n555), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1340gat));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n205), .A3(new_n633), .ZN(new_n839));
  OAI21_X1  g638(.A(G120gat), .B1(new_n834), .B2(new_n634), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1341gat));
  NOR2_X1   g640(.A1(new_n834), .A2(new_n658), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(new_n209), .ZN(G1342gat));
  OR2_X1    g642(.A1(new_n834), .A2(new_n607), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .A3(new_n214), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(G134gat), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT56), .B1(new_n844), .B2(new_n214), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  NOR3_X1   g647(.A1(new_n652), .A2(new_n639), .A3(new_n424), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n555), .A2(new_n801), .A3(new_n823), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n816), .B(KEYINPUT118), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n607), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n574), .B1(new_n853), .B2(new_n825), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n680), .B1(new_n854), .B2(new_n793), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n850), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n829), .A2(new_n857), .A3(new_n680), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n229), .B1(new_n859), .B2(new_n554), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n808), .A2(KEYINPUT115), .A3(new_n816), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n808), .B2(new_n816), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n861), .A2(new_n862), .A3(new_n606), .ZN(new_n863));
  INV_X1    g662(.A(new_n825), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n658), .A3(new_n826), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n419), .B1(new_n866), .B2(new_n794), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n849), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G141gat), .A3(new_n555), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT58), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n555), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n858), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT119), .A4(new_n871), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n874), .A2(G141gat), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n869), .A2(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(new_n868), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n227), .A3(new_n633), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  AOI211_X1 g682(.A(KEYINPUT59), .B(new_n227), .C1(new_n859), .C2(new_n633), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n829), .A2(new_n680), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n635), .A2(new_n871), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n857), .B(new_n680), .C1(new_n854), .C2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n887), .A2(new_n633), .A3(new_n849), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n882), .A2(new_n883), .B1(new_n884), .B2(new_n891), .ZN(G1345gat));
  NAND4_X1  g691(.A1(new_n859), .A2(new_n234), .A3(new_n235), .A4(new_n574), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n868), .A2(new_n658), .B1(new_n249), .B2(new_n248), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1346gat));
  NAND2_X1  g694(.A1(new_n859), .A2(new_n606), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n859), .A2(KEYINPUT121), .A3(new_n606), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(G162gat), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n222), .A3(new_n606), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n640), .A2(new_n488), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n832), .B(new_n904), .C1(new_n866), .C2(new_n794), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n555), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n300), .A3(new_n554), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1348gat));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n633), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g710(.A1(new_n905), .A2(new_n574), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G183gat), .ZN(new_n913));
  INV_X1    g712(.A(new_n316), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n912), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT60), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  OAI221_X1 g717(.A(new_n913), .B1(KEYINPUT122), .B2(new_n918), .C1(new_n914), .C2(new_n912), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1350gat));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n922), .A3(new_n314), .A4(new_n606), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n829), .A2(new_n831), .A3(new_n606), .A4(new_n903), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n924), .B2(G190gat), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(G190gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(KEYINPUT61), .A3(G190gat), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n921), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n923), .A2(new_n925), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n933), .A2(KEYINPUT124), .A3(new_n930), .A4(new_n929), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n904), .A2(new_n652), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n889), .B(new_n936), .C1(new_n867), .C2(new_n857), .ZN(new_n937));
  OAI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n555), .ZN(new_n938));
  INV_X1    g737(.A(new_n936), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n886), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(G197gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n554), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n942), .ZN(G1352gat));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n617), .A3(new_n633), .ZN(new_n944));
  AND2_X1   g743(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n945));
  NOR2_X1   g744(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n887), .A2(new_n633), .A3(new_n889), .ZN(new_n948));
  OAI21_X1  g747(.A(G204gat), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n947), .B(new_n949), .C1(new_n945), .C2(new_n944), .ZN(G1353gat));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g752(.A(G211gat), .B(new_n953), .C1(new_n937), .C2(new_n658), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n352), .A3(new_n574), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n955), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G1354gat));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n937), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n606), .B1(new_n937), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g761(.A(G218gat), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n940), .A2(new_n353), .A3(new_n606), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


