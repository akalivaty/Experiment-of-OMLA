

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786;

  XNOR2_X1 U379 ( .A(G143), .B(G104), .ZN(n504) );
  XNOR2_X1 U380 ( .A(G101), .B(G107), .ZN(n463) );
  INV_X2 U381 ( .A(n382), .ZN(n383) );
  XNOR2_X2 U382 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  XNOR2_X2 U383 ( .A(n358), .B(n657), .ZN(n659) );
  XNOR2_X2 U384 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X2 U385 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X2 U386 ( .A(n651), .B(KEYINPUT122), .ZN(n652) );
  NAND2_X2 U387 ( .A1(n414), .A2(n366), .ZN(n586) );
  XNOR2_X1 U388 ( .A(KEYINPUT18), .B(KEYINPUT93), .ZN(n481) );
  XOR2_X1 U389 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n498) );
  XOR2_X1 U390 ( .A(G140), .B(G122), .Z(n503) );
  INV_X1 U391 ( .A(G237), .ZN(n437) );
  INV_X1 U392 ( .A(G137), .ZN(n452) );
  XOR2_X1 U393 ( .A(n360), .B(n403), .Z(n356) );
  AND2_X2 U394 ( .A1(n408), .A2(n406), .ZN(n412) );
  XNOR2_X2 U395 ( .A(n357), .B(n463), .ZN(n777) );
  NAND2_X2 U396 ( .A1(n393), .A2(n392), .ZN(n621) );
  AND2_X2 U397 ( .A1(n398), .A2(n363), .ZN(n393) );
  AND2_X4 U398 ( .A1(n650), .A2(n649), .ZN(n743) );
  OR2_X2 U399 ( .A1(n745), .A2(G902), .ZN(n470) );
  OR2_X1 U400 ( .A1(n579), .A2(n708), .ZN(n537) );
  OR2_X1 U401 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X2 U402 ( .A(n777), .B(KEYINPUT66), .ZN(n488) );
  XNOR2_X2 U403 ( .A(n517), .B(n427), .ZN(n727) );
  XNOR2_X2 U404 ( .A(n480), .B(G134), .ZN(n517) );
  NOR2_X2 U405 ( .A1(n642), .A2(n643), .ZN(n638) );
  XNOR2_X1 U406 ( .A(n468), .B(n435), .ZN(n658) );
  AND2_X1 U407 ( .A1(n410), .A2(n584), .ZN(n409) );
  AND2_X1 U408 ( .A1(n414), .A2(KEYINPUT84), .ZN(n407) );
  NAND2_X1 U409 ( .A1(n370), .A2(KEYINPUT82), .ZN(n414) );
  NOR2_X1 U410 ( .A1(n720), .A2(n619), .ZN(n610) );
  XNOR2_X1 U411 ( .A(G104), .B(KEYINPUT70), .ZN(n464) );
  NAND2_X1 U412 ( .A1(n374), .A2(n371), .ZN(n378) );
  AND2_X1 U413 ( .A1(n376), .A2(n364), .ZN(n374) );
  NAND2_X1 U414 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U415 ( .A1(n404), .A2(n590), .ZN(n411) );
  AND2_X1 U416 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X1 U417 ( .A1(n585), .A2(n587), .ZN(n410) );
  NAND2_X1 U418 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U419 ( .A1(n554), .A2(n569), .ZN(n555) );
  XNOR2_X1 U420 ( .A(n571), .B(n570), .ZN(n719) );
  XNOR2_X1 U421 ( .A(n458), .B(n457), .ZN(n558) );
  XNOR2_X1 U422 ( .A(n545), .B(KEYINPUT6), .ZN(n563) );
  BUF_X1 U423 ( .A(n658), .Z(n358) );
  NAND2_X1 U424 ( .A1(n780), .A2(G234), .ZN(n449) );
  XNOR2_X1 U425 ( .A(n464), .B(G110), .ZN(n357) );
  XNOR2_X2 U426 ( .A(G101), .B(G116), .ZN(n429) );
  XNOR2_X1 U427 ( .A(KEYINPUT72), .B(KEYINPUT65), .ZN(n443) );
  XNOR2_X2 U428 ( .A(G137), .B(KEYINPUT5), .ZN(n428) );
  XNOR2_X2 U429 ( .A(G146), .B(G125), .ZN(n478) );
  NAND2_X1 U430 ( .A1(n584), .A2(n585), .ZN(n405) );
  BUF_X1 U431 ( .A(n777), .Z(n359) );
  NAND2_X1 U432 ( .A1(n393), .A2(n392), .ZN(n360) );
  XNOR2_X1 U433 ( .A(n621), .B(n403), .ZN(n532) );
  XNOR2_X1 U434 ( .A(n396), .B(n576), .ZN(n593) );
  BUF_X1 U435 ( .A(n593), .Z(n726) );
  NAND2_X1 U436 ( .A1(n593), .A2(KEYINPUT44), .ZN(n585) );
  NAND2_X1 U437 ( .A1(n477), .A2(G224), .ZN(n390) );
  XNOR2_X1 U438 ( .A(n369), .B(KEYINPUT77), .ZN(n368) );
  NAND2_X1 U439 ( .A1(n380), .A2(n379), .ZN(n369) );
  XNOR2_X2 U440 ( .A(n544), .B(n365), .ZN(n554) );
  XNOR2_X1 U441 ( .A(n592), .B(KEYINPUT85), .ZN(n597) );
  NAND2_X1 U442 ( .A1(n412), .A2(n411), .ZN(n591) );
  NOR2_X1 U443 ( .A1(n420), .A2(KEYINPUT82), .ZN(n419) );
  INV_X2 U444 ( .A(G953), .ZN(n477) );
  INV_X1 U445 ( .A(KEYINPUT101), .ZN(n415) );
  INV_X1 U446 ( .A(n641), .ZN(n379) );
  INV_X1 U447 ( .A(KEYINPUT12), .ZN(n384) );
  XNOR2_X1 U448 ( .A(G113), .B(G131), .ZN(n502) );
  XNOR2_X1 U449 ( .A(KEYINPUT4), .B(G131), .ZN(n427) );
  AND2_X1 U450 ( .A1(n563), .A2(n568), .ZN(n423) );
  NOR2_X1 U451 ( .A1(n648), .A2(n381), .ZN(n682) );
  INV_X1 U452 ( .A(G902), .ZN(n520) );
  XNOR2_X1 U453 ( .A(n638), .B(KEYINPUT79), .ZN(n730) );
  NAND2_X1 U454 ( .A1(n425), .A2(n426), .ZN(n614) );
  INV_X1 U455 ( .A(KEYINPUT19), .ZN(n403) );
  NOR2_X1 U456 ( .A1(n418), .A2(n417), .ZN(n416) );
  NOR2_X1 U457 ( .A1(n697), .A2(n556), .ZN(n418) );
  INV_X1 U458 ( .A(n421), .ZN(n370) );
  INV_X1 U459 ( .A(KEYINPUT119), .ZN(n372) );
  OR2_X1 U460 ( .A1(n723), .A2(KEYINPUT119), .ZN(n375) );
  XNOR2_X1 U461 ( .A(n553), .B(n401), .ZN(n400) );
  INV_X1 U462 ( .A(KEYINPUT64), .ZN(n401) );
  INV_X1 U463 ( .A(n700), .ZN(n417) );
  AND2_X1 U464 ( .A1(n527), .A2(KEYINPUT86), .ZN(n361) );
  AND2_X1 U465 ( .A1(n531), .A2(n530), .ZN(n362) );
  OR2_X1 U466 ( .A1(n527), .A2(KEYINPUT86), .ZN(n363) );
  AND2_X1 U467 ( .A1(n375), .A2(n780), .ZN(n364) );
  XOR2_X1 U468 ( .A(n543), .B(KEYINPUT22), .Z(n365) );
  INV_X1 U469 ( .A(KEYINPUT82), .ZN(n556) );
  INV_X1 U470 ( .A(n568), .ZN(n696) );
  XNOR2_X2 U471 ( .A(n436), .B(G472), .ZN(n545) );
  XNOR2_X2 U472 ( .A(n727), .B(G146), .ZN(n468) );
  NAND2_X1 U473 ( .A1(n407), .A2(n366), .ZN(n406) );
  AND2_X2 U474 ( .A1(n413), .A2(n416), .ZN(n366) );
  NAND2_X1 U475 ( .A1(n367), .A2(n424), .ZN(n650) );
  NAND2_X1 U476 ( .A1(n368), .A2(n639), .ZN(n367) );
  XNOR2_X2 U477 ( .A(n555), .B(KEYINPUT81), .ZN(n421) );
  INV_X1 U478 ( .A(n724), .ZN(n373) );
  NAND2_X1 U479 ( .A1(n724), .A2(n377), .ZN(n376) );
  AND2_X1 U480 ( .A1(n723), .A2(KEYINPUT119), .ZN(n377) );
  XNOR2_X1 U481 ( .A(n378), .B(n725), .ZN(G75) );
  XNOR2_X1 U482 ( .A(n602), .B(KEYINPUT45), .ZN(n380) );
  XNOR2_X2 U483 ( .A(G116), .B(G122), .ZN(n515) );
  XNOR2_X1 U484 ( .A(n602), .B(n601), .ZN(n381) );
  INV_X1 U485 ( .A(n743), .ZN(n382) );
  XNOR2_X1 U486 ( .A(n499), .B(n384), .ZN(n501) );
  XNOR2_X1 U487 ( .A(n395), .B(n415), .ZN(n394) );
  NAND2_X1 U488 ( .A1(n397), .A2(n574), .ZN(n396) );
  NAND2_X1 U489 ( .A1(n483), .A2(n482), .ZN(n387) );
  NAND2_X1 U490 ( .A1(n385), .A2(n386), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n388), .A2(n387), .ZN(n486) );
  INV_X1 U492 ( .A(n483), .ZN(n385) );
  INV_X1 U493 ( .A(n482), .ZN(n386) );
  XNOR2_X1 U494 ( .A(n389), .B(KEYINPUT34), .ZN(n397) );
  NOR2_X1 U495 ( .A1(n579), .A2(n719), .ZN(n389) );
  XNOR2_X1 U496 ( .A(n391), .B(n390), .ZN(n479) );
  XNOR2_X2 U497 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n391) );
  NAND2_X1 U498 ( .A1(n532), .A2(n362), .ZN(n533) );
  NAND2_X1 U499 ( .A1(n399), .A2(n529), .ZN(n392) );
  NAND2_X1 U500 ( .A1(n394), .A2(n583), .ZN(n584) );
  NAND2_X1 U501 ( .A1(n765), .A2(n752), .ZN(n395) );
  XNOR2_X2 U502 ( .A(n581), .B(n580), .ZN(n752) );
  XNOR2_X2 U503 ( .A(n537), .B(n536), .ZN(n765) );
  NAND2_X1 U504 ( .A1(n528), .A2(n361), .ZN(n398) );
  XNOR2_X2 U505 ( .A(n422), .B(n492), .ZN(n528) );
  INV_X1 U506 ( .A(n528), .ZN(n399) );
  NAND2_X1 U507 ( .A1(n400), .A2(n417), .ZN(n588) );
  XNOR2_X2 U508 ( .A(n402), .B(KEYINPUT32), .ZN(n589) );
  NAND2_X1 U509 ( .A1(n549), .A2(n548), .ZN(n402) );
  NOR2_X2 U510 ( .A1(n772), .A2(G237), .ZN(n496) );
  NAND2_X1 U511 ( .A1(n405), .A2(KEYINPUT84), .ZN(n404) );
  NAND2_X1 U512 ( .A1(n409), .A2(n586), .ZN(n408) );
  NAND2_X1 U513 ( .A1(n421), .A2(n419), .ZN(n413) );
  INV_X1 U514 ( .A(n697), .ZN(n420) );
  NAND2_X1 U515 ( .A1(n665), .A2(n641), .ZN(n422) );
  XNOR2_X1 U516 ( .A(n487), .B(n488), .ZN(n665) );
  INV_X1 U517 ( .A(n563), .ZN(n569) );
  NAND2_X1 U518 ( .A1(n625), .A2(n423), .ZN(n571) );
  OR2_X1 U519 ( .A1(n641), .A2(n640), .ZN(n424) );
  XNOR2_X1 U520 ( .A(KEYINPUT30), .B(n440), .ZN(n425) );
  XOR2_X1 U521 ( .A(n476), .B(KEYINPUT71), .Z(n426) );
  INV_X1 U522 ( .A(n786), .ZN(n611) );
  XNOR2_X1 U523 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U524 ( .A(n431), .B(n430), .ZN(n434) );
  INV_X1 U525 ( .A(n730), .ZN(n639) );
  INV_X1 U526 ( .A(KEYINPUT78), .ZN(n684) );
  INV_X1 U527 ( .A(n682), .ZN(n649) );
  XNOR2_X2 U528 ( .A(G143), .B(G128), .ZN(n480) );
  BUF_X2 U529 ( .A(G953), .Z(n772) );
  NAND2_X1 U530 ( .A1(n496), .A2(G210), .ZN(n430) );
  XNOR2_X1 U531 ( .A(G119), .B(G113), .ZN(n433) );
  XNOR2_X1 U532 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X1 U533 ( .A(n433), .B(n432), .ZN(n485) );
  XNOR2_X1 U534 ( .A(n434), .B(n485), .ZN(n435) );
  NOR2_X2 U535 ( .A1(n658), .A2(G902), .ZN(n436) );
  XNOR2_X1 U536 ( .A(n545), .B(KEYINPUT107), .ZN(n606) );
  INV_X1 U537 ( .A(n606), .ZN(n551) );
  NAND2_X1 U538 ( .A1(n520), .A2(n437), .ZN(n489) );
  NAND2_X1 U539 ( .A1(n489), .A2(G214), .ZN(n439) );
  INV_X1 U540 ( .A(KEYINPUT96), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n439), .B(n438), .ZN(n686) );
  NOR2_X1 U542 ( .A1(n551), .A2(n686), .ZN(n440) );
  XOR2_X1 U543 ( .A(KEYINPUT24), .B(G110), .Z(n442) );
  XNOR2_X1 U544 ( .A(G119), .B(G128), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n442), .B(n441), .ZN(n447) );
  INV_X1 U546 ( .A(n443), .ZN(n445) );
  XNOR2_X1 U547 ( .A(KEYINPUT76), .B(KEYINPUT23), .ZN(n444) );
  XNOR2_X1 U548 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U549 ( .A(n447), .B(n446), .ZN(n448) );
  INV_X1 U550 ( .A(n448), .ZN(n451) );
  BUF_X4 U551 ( .A(n477), .Z(n780) );
  XOR2_X1 U552 ( .A(KEYINPUT8), .B(n449), .Z(n511) );
  NAND2_X1 U553 ( .A1(n511), .A2(G221), .ZN(n450) );
  XNOR2_X1 U554 ( .A(n451), .B(n450), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n478), .B(KEYINPUT10), .ZN(n500) );
  XNOR2_X1 U556 ( .A(n452), .B(G140), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n500), .B(n466), .ZN(n728) );
  XNOR2_X1 U558 ( .A(n453), .B(n728), .ZN(n651) );
  NAND2_X1 U559 ( .A1(n651), .A2(n520), .ZN(n458) );
  XOR2_X1 U560 ( .A(KEYINPUT20), .B(KEYINPUT97), .Z(n455) );
  NAND2_X1 U561 ( .A1(G234), .A2(n641), .ZN(n454) );
  XNOR2_X1 U562 ( .A(n455), .B(n454), .ZN(n459) );
  NAND2_X1 U563 ( .A1(n459), .A2(G217), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n459), .A2(G221), .ZN(n461) );
  INV_X1 U566 ( .A(KEYINPUT21), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n699) );
  INV_X1 U568 ( .A(KEYINPUT98), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n699), .B(n462), .ZN(n541) );
  NOR2_X2 U570 ( .A1(n558), .A2(n541), .ZN(n568) );
  NAND2_X1 U571 ( .A1(n780), .A2(G227), .ZN(n465) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n488), .B(n467), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n469), .B(n468), .ZN(n745) );
  XNOR2_X2 U575 ( .A(n470), .B(G469), .ZN(n608) );
  NAND2_X1 U576 ( .A1(n568), .A2(n608), .ZN(n577) );
  NAND2_X1 U577 ( .A1(G234), .A2(G237), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n471), .B(KEYINPUT14), .ZN(n716) );
  INV_X1 U579 ( .A(G952), .ZN(n654) );
  NAND2_X1 U580 ( .A1(n780), .A2(n654), .ZN(n473) );
  NAND2_X1 U581 ( .A1(n772), .A2(n520), .ZN(n472) );
  AND2_X1 U582 ( .A1(n473), .A2(n472), .ZN(n474) );
  AND2_X1 U583 ( .A1(n716), .A2(n474), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n772), .A2(G900), .ZN(n475) );
  NAND2_X1 U585 ( .A1(n531), .A2(n475), .ZN(n559) );
  NOR2_X1 U586 ( .A1(n577), .A2(n559), .ZN(n476) );
  XNOR2_X1 U587 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U588 ( .A(n480), .B(n481), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n515), .B(KEYINPUT16), .ZN(n484) );
  XNOR2_X1 U590 ( .A(n485), .B(n484), .ZN(n778) );
  XNOR2_X1 U591 ( .A(n486), .B(n778), .ZN(n487) );
  NAND2_X1 U592 ( .A1(n489), .A2(G210), .ZN(n491) );
  XNOR2_X1 U593 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n492) );
  BUF_X1 U595 ( .A(n528), .Z(n493) );
  XNOR2_X1 U596 ( .A(n493), .B(KEYINPUT38), .ZN(n687) );
  NOR2_X1 U597 ( .A1(n614), .A2(n687), .ZN(n495) );
  XNOR2_X1 U598 ( .A(KEYINPUT80), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U599 ( .A(n495), .B(n494), .ZN(n524) );
  XNOR2_X1 U600 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n509) );
  NAND2_X1 U601 ( .A1(G214), .A2(n496), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U603 ( .A(n501), .B(n500), .ZN(n507) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n507), .B(n506), .ZN(n675) );
  NOR2_X1 U607 ( .A1(G902), .A2(n675), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U609 ( .A(n510), .B(G475), .ZN(n573) );
  XOR2_X1 U610 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n513) );
  NAND2_X1 U611 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n513), .B(n512), .ZN(n519) );
  XNOR2_X1 U613 ( .A(G107), .B(KEYINPUT9), .ZN(n514) );
  XNOR2_X1 U614 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U615 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U616 ( .A(n519), .B(n518), .ZN(n738) );
  NAND2_X1 U617 ( .A1(n738), .A2(n520), .ZN(n521) );
  XNOR2_X1 U618 ( .A(n521), .B(G478), .ZN(n540) );
  NAND2_X1 U619 ( .A1(n573), .A2(n540), .ZN(n522) );
  XNOR2_X1 U620 ( .A(n522), .B(KEYINPUT105), .ZN(n757) );
  INV_X1 U621 ( .A(KEYINPUT106), .ZN(n523) );
  XNOR2_X1 U622 ( .A(n757), .B(n523), .ZN(n582) );
  NOR2_X1 U623 ( .A1(n524), .A2(n582), .ZN(n643) );
  XOR2_X1 U624 ( .A(G134), .B(n643), .Z(G36) );
  OR2_X1 U625 ( .A1(n573), .A2(n540), .ZN(n764) );
  NOR2_X1 U626 ( .A1(n524), .A2(n764), .ZN(n526) );
  XNOR2_X1 U627 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n603) );
  XOR2_X1 U629 ( .A(G131), .B(n603), .Z(G33) );
  INV_X1 U630 ( .A(n686), .ZN(n527) );
  INV_X1 U631 ( .A(KEYINPUT86), .ZN(n529) );
  NAND2_X1 U632 ( .A1(n772), .A2(G898), .ZN(n530) );
  XNOR2_X2 U633 ( .A(n533), .B(KEYINPUT0), .ZN(n579) );
  XNOR2_X2 U634 ( .A(n608), .B(KEYINPUT1), .ZN(n625) );
  INV_X1 U635 ( .A(n625), .ZN(n550) );
  INV_X1 U636 ( .A(n545), .ZN(n704) );
  NAND2_X1 U637 ( .A1(n568), .A2(n704), .ZN(n534) );
  OR2_X1 U638 ( .A1(n550), .A2(n534), .ZN(n708) );
  INV_X1 U639 ( .A(KEYINPUT100), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n535), .B(KEYINPUT31), .ZN(n536) );
  INV_X1 U641 ( .A(n765), .ZN(n538) );
  NAND2_X1 U642 ( .A1(n538), .A2(n757), .ZN(n539) );
  XNOR2_X1 U643 ( .A(n539), .B(G116), .ZN(G18) );
  INV_X1 U644 ( .A(n540), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n689) );
  OR2_X1 U646 ( .A1(n689), .A2(n541), .ZN(n542) );
  NOR2_X2 U647 ( .A1(n579), .A2(n542), .ZN(n544) );
  INV_X1 U648 ( .A(KEYINPUT68), .ZN(n543) );
  BUF_X1 U649 ( .A(n554), .Z(n549) );
  XNOR2_X1 U650 ( .A(n569), .B(KEYINPUT74), .ZN(n547) );
  AND2_X1 U651 ( .A1(n625), .A2(n558), .ZN(n546) );
  AND2_X1 U652 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U653 ( .A(n589), .B(G119), .ZN(G21) );
  BUF_X1 U654 ( .A(n550), .Z(n697) );
  AND2_X1 U655 ( .A1(n697), .A2(n551), .ZN(n552) );
  NAND2_X1 U656 ( .A1(n554), .A2(n552), .ZN(n553) );
  INV_X1 U657 ( .A(n558), .ZN(n700) );
  XNOR2_X1 U658 ( .A(n588), .B(G110), .ZN(G12) );
  BUF_X1 U659 ( .A(n586), .Z(n557) );
  XNOR2_X1 U660 ( .A(n557), .B(G101), .ZN(G3) );
  NAND2_X1 U661 ( .A1(n558), .A2(n699), .ZN(n560) );
  NOR2_X1 U662 ( .A1(n560), .A2(n559), .ZN(n605) );
  INV_X1 U663 ( .A(n605), .ZN(n561) );
  NOR2_X1 U664 ( .A1(n764), .A2(n561), .ZN(n562) );
  NAND2_X1 U665 ( .A1(n563), .A2(n562), .ZN(n623) );
  NOR2_X1 U666 ( .A1(n686), .A2(n623), .ZN(n564) );
  XNOR2_X1 U667 ( .A(KEYINPUT108), .B(n564), .ZN(n565) );
  NAND2_X1 U668 ( .A1(n565), .A2(n697), .ZN(n566) );
  XNOR2_X1 U669 ( .A(n566), .B(KEYINPUT43), .ZN(n567) );
  NAND2_X1 U670 ( .A1(n567), .A2(n399), .ZN(n636) );
  XNOR2_X1 U671 ( .A(n636), .B(G140), .ZN(G42) );
  XNOR2_X1 U672 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n570) );
  OR2_X1 U673 ( .A1(n573), .A2(n572), .ZN(n617) );
  INV_X1 U674 ( .A(n617), .ZN(n574) );
  INV_X1 U675 ( .A(KEYINPUT73), .ZN(n575) );
  XNOR2_X1 U676 ( .A(n575), .B(KEYINPUT35), .ZN(n576) );
  OR2_X1 U677 ( .A1(n577), .A2(n704), .ZN(n578) );
  INV_X1 U678 ( .A(KEYINPUT99), .ZN(n580) );
  AND2_X1 U679 ( .A1(n582), .A2(n764), .ZN(n691) );
  INV_X1 U680 ( .A(n691), .ZN(n583) );
  INV_X1 U681 ( .A(KEYINPUT84), .ZN(n587) );
  NAND2_X1 U682 ( .A1(n592), .A2(KEYINPUT44), .ZN(n590) );
  XNOR2_X1 U683 ( .A(n591), .B(KEYINPUT83), .ZN(n600) );
  INV_X1 U684 ( .A(n726), .ZN(n595) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n594) );
  AND2_X1 U686 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U687 ( .A(n598), .B(KEYINPUT67), .ZN(n599) );
  NAND2_X1 U688 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U689 ( .A(KEYINPUT45), .ZN(n601) );
  INV_X1 U690 ( .A(n603), .ZN(n612) );
  OR2_X1 U691 ( .A1(n687), .A2(n686), .ZN(n690) );
  NOR2_X1 U692 ( .A1(n689), .A2(n690), .ZN(n604) );
  XNOR2_X1 U693 ( .A(KEYINPUT41), .B(n604), .ZN(n720) );
  NAND2_X1 U694 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U695 ( .A(KEYINPUT28), .B(n607), .Z(n609) );
  NAND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n610), .B(KEYINPUT42), .ZN(n786) );
  NAND2_X1 U698 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U699 ( .A(n613), .B(KEYINPUT46), .ZN(n634) );
  INV_X1 U700 ( .A(n614), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n615), .A2(n493), .ZN(n616) );
  XOR2_X1 U702 ( .A(KEYINPUT109), .B(n616), .Z(n618) );
  NOR2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n760) );
  AND2_X1 U704 ( .A1(n691), .A2(KEYINPUT69), .ZN(n620) );
  NOR2_X1 U705 ( .A1(n619), .A2(n356), .ZN(n762) );
  NAND2_X1 U706 ( .A1(n620), .A2(n762), .ZN(n627) );
  INV_X1 U707 ( .A(n360), .ZN(n622) );
  NOR2_X1 U708 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U709 ( .A(n624), .B(KEYINPUT36), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n626), .A2(n420), .ZN(n769) );
  NAND2_X1 U711 ( .A1(n627), .A2(n769), .ZN(n628) );
  NOR2_X1 U712 ( .A1(n760), .A2(n628), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n691), .A2(KEYINPUT69), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n629), .A2(n762), .ZN(n630) );
  XOR2_X1 U715 ( .A(KEYINPUT47), .B(n630), .Z(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U718 ( .A(n635), .B(KEYINPUT48), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n642) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n640) );
  INV_X1 U721 ( .A(n642), .ZN(n647) );
  INV_X1 U722 ( .A(n643), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(KEYINPUT75), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n743), .A2(G217), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n654), .A2(n772), .ZN(n741) );
  NAND2_X1 U729 ( .A1(n655), .A2(n741), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U731 ( .A1(n743), .A2(G472), .ZN(n660) );
  XNOR2_X1 U732 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n661), .A2(n741), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT87), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G57) );
  NAND2_X1 U738 ( .A1(n743), .A2(G210), .ZN(n670) );
  BUF_X1 U739 ( .A(n665), .Z(n668) );
  XNOR2_X1 U740 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n666) );
  XOR2_X1 U741 ( .A(n666), .B(KEYINPUT55), .Z(n667) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(n741), .ZN(n673) );
  XOR2_X1 U744 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(G51) );
  NAND2_X1 U746 ( .A1(n743), .A2(G475), .ZN(n677) );
  XNOR2_X1 U747 ( .A(KEYINPUT90), .B(KEYINPUT59), .ZN(n674) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n678), .A2(n741), .ZN(n680) );
  INV_X1 U750 ( .A(KEYINPUT60), .ZN(n679) );
  XNOR2_X1 U751 ( .A(n680), .B(n679), .ZN(G60) );
  NOR2_X1 U752 ( .A1(n730), .A2(n381), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n681), .A2(KEYINPUT2), .ZN(n683) );
  NOR2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(n724) );
  AND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT118), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n695), .A2(n719), .ZN(n714) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n698), .B(KEYINPUT50), .ZN(n707) );
  XOR2_X1 U764 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n702) );
  OR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U766 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U767 ( .A(n703), .B(KEYINPUT116), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n710) );
  XNOR2_X1 U772 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U773 ( .A1(n712), .A2(n720), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n715), .B(KEYINPUT52), .ZN(n718) );
  NAND2_X1 U776 ( .A1(G952), .A2(n716), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n722), .A2(n721), .ZN(n723) );
  INV_X1 U780 ( .A(KEYINPUT53), .ZN(n725) );
  XOR2_X1 U781 ( .A(n726), .B(G122), .Z(G24) );
  XNOR2_X1 U782 ( .A(n727), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n730), .B(n732), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n731), .A2(n780), .ZN(n737) );
  XOR2_X1 U786 ( .A(n732), .B(KEYINPUT127), .Z(n733) );
  XNOR2_X1 U787 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U788 ( .A1(G900), .A2(n734), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n735), .A2(n772), .ZN(n736) );
  NAND2_X1 U790 ( .A1(n737), .A2(n736), .ZN(G72) );
  NAND2_X1 U791 ( .A1(n383), .A2(G478), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n738), .B(KEYINPUT121), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n742) );
  INV_X1 U794 ( .A(n741), .ZN(n748) );
  NOR2_X1 U795 ( .A1(n742), .A2(n748), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n383), .A2(G469), .ZN(n747) );
  XOR2_X1 U797 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n747), .B(n746), .ZN(n749) );
  NOR2_X1 U800 ( .A1(n749), .A2(n748), .ZN(G54) );
  NOR2_X1 U801 ( .A1(n752), .A2(n764), .ZN(n750) );
  XOR2_X1 U802 ( .A(KEYINPUT112), .B(n750), .Z(n751) );
  XNOR2_X1 U803 ( .A(G104), .B(n751), .ZN(G6) );
  INV_X1 U804 ( .A(n752), .ZN(n753) );
  NAND2_X1 U805 ( .A1(n753), .A2(n757), .ZN(n755) );
  XOR2_X1 U806 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n754) );
  XNOR2_X1 U807 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U808 ( .A(G107), .B(n756), .ZN(G9) );
  XOR2_X1 U809 ( .A(G128), .B(KEYINPUT29), .Z(n759) );
  NAND2_X1 U810 ( .A1(n762), .A2(n757), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n759), .B(n758), .ZN(G30) );
  XOR2_X1 U812 ( .A(G143), .B(n760), .Z(G45) );
  INV_X1 U813 ( .A(n764), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(G146), .ZN(G48) );
  XOR2_X1 U816 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n767) );
  NOR2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U818 ( .A(n767), .B(n766), .Z(n768) );
  XNOR2_X1 U819 ( .A(G113), .B(n768), .ZN(G15) );
  XOR2_X1 U820 ( .A(G125), .B(n769), .Z(n770) );
  XNOR2_X1 U821 ( .A(n770), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U822 ( .A(n381), .ZN(n771) );
  NAND2_X1 U823 ( .A1(n771), .A2(n780), .ZN(n776) );
  NAND2_X1 U824 ( .A1(n772), .A2(G224), .ZN(n773) );
  XNOR2_X1 U825 ( .A(KEYINPUT61), .B(n773), .ZN(n774) );
  NAND2_X1 U826 ( .A1(n774), .A2(G898), .ZN(n775) );
  NAND2_X1 U827 ( .A1(n776), .A2(n775), .ZN(n784) );
  XNOR2_X1 U828 ( .A(n359), .B(KEYINPUT124), .ZN(n779) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(n782) );
  NOR2_X1 U830 ( .A1(n780), .A2(G898), .ZN(n781) );
  NOR2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U832 ( .A(n784), .B(n783), .ZN(n785) );
  XOR2_X1 U833 ( .A(KEYINPUT125), .B(n785), .Z(G69) );
  XOR2_X1 U834 ( .A(G137), .B(n786), .Z(G39) );
endmodule

