

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n751, n752, n753, n754, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792;

  AND2_X1 U370 ( .A1(n358), .A2(n357), .ZN(n751) );
  AND2_X1 U371 ( .A1(n361), .A2(n360), .ZN(n756) );
  AND2_X1 U372 ( .A1(n364), .A2(n363), .ZN(n680) );
  INV_X1 U373 ( .A(n762), .ZN(n357) );
  INV_X1 U374 ( .A(n762), .ZN(n360) );
  INV_X1 U375 ( .A(n762), .ZN(n363) );
  BUF_X1 U376 ( .A(n737), .Z(n352) );
  XNOR2_X1 U377 ( .A(n614), .B(KEYINPUT46), .ZN(n615) );
  NAND2_X1 U378 ( .A1(n413), .A2(n410), .ZN(n419) );
  NAND2_X1 U379 ( .A1(n440), .A2(n439), .ZN(n504) );
  NAND2_X1 U380 ( .A1(n438), .A2(n437), .ZN(n792) );
  BUF_X1 U381 ( .A(n710), .Z(n351) );
  XNOR2_X1 U382 ( .A(n356), .B(n648), .ZN(n654) );
  INV_X1 U383 ( .A(n447), .ZN(n353) );
  XNOR2_X1 U384 ( .A(n403), .B(n594), .ZN(n710) );
  XNOR2_X1 U385 ( .A(n601), .B(KEYINPUT38), .ZN(n724) );
  INV_X1 U386 ( .A(n625), .ZN(n601) );
  XNOR2_X1 U387 ( .A(n593), .B(n592), .ZN(n403) );
  NOR2_X1 U388 ( .A1(G902), .A2(n668), .ZN(n593) );
  INV_X1 U389 ( .A(n712), .ZN(n660) );
  XNOR2_X1 U390 ( .A(KEYINPUT71), .B(G472), .ZN(n584) );
  XOR2_X1 U391 ( .A(n397), .B(n435), .Z(n368) );
  XNOR2_X1 U392 ( .A(n514), .B(n513), .ZN(n576) );
  XNOR2_X1 U393 ( .A(G119), .B(G113), .ZN(n513) );
  BUF_X1 U394 ( .A(n673), .Z(n350) );
  NOR2_X2 U395 ( .A1(G952), .A2(n531), .ZN(n762) );
  NOR2_X1 U396 ( .A1(n354), .A2(n353), .ZN(n438) );
  INV_X1 U397 ( .A(n448), .ZN(n354) );
  NAND2_X1 U398 ( .A1(n759), .A2(G217), .ZN(n760) );
  AND2_X4 U399 ( .A1(n454), .A2(n460), .ZN(n759) );
  NOR2_X2 U400 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U401 ( .A1(n355), .A2(n449), .ZN(n747) );
  NAND2_X1 U402 ( .A1(n452), .A2(n453), .ZN(n355) );
  NOR2_X2 U403 ( .A1(n646), .A2(n491), .ZN(n356) );
  AND2_X2 U404 ( .A1(n463), .A2(n402), .ZN(n658) );
  XNOR2_X1 U405 ( .A(n748), .B(n359), .ZN(n358) );
  INV_X1 U406 ( .A(n749), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n753), .B(n362), .ZN(n361) );
  INV_X1 U408 ( .A(n754), .ZN(n362) );
  XNOR2_X1 U409 ( .A(n676), .B(n365), .ZN(n364) );
  INV_X1 U410 ( .A(n677), .ZN(n365) );
  XNOR2_X1 U411 ( .A(G122), .B(G113), .ZN(n540) );
  INV_X1 U412 ( .A(G953), .ZN(n531) );
  AND2_X2 U413 ( .A1(n458), .A2(n380), .ZN(n456) );
  XNOR2_X2 U414 ( .A(n637), .B(n636), .ZN(n646) );
  NOR2_X2 U415 ( .A1(n428), .A2(n635), .ZN(n637) );
  NOR2_X1 U416 ( .A1(n620), .A2(n724), .ZN(n478) );
  AND2_X1 U417 ( .A1(n406), .A2(n407), .ZN(n405) );
  NOR2_X1 U418 ( .A1(n382), .A2(n790), .ZN(n482) );
  AND2_X1 U419 ( .A1(n417), .A2(n414), .ZN(n413) );
  XNOR2_X1 U420 ( .A(n367), .B(KEYINPUT110), .ZN(n790) );
  XNOR2_X1 U421 ( .A(n478), .B(n613), .ZN(n629) );
  AND2_X1 U422 ( .A1(n598), .A2(n601), .ZN(n599) );
  NOR2_X1 U423 ( .A1(n586), .A2(n469), .ZN(n598) );
  XNOR2_X1 U424 ( .A(n585), .B(KEYINPUT103), .ZN(n586) );
  NOR2_X1 U425 ( .A1(n650), .A2(n603), .ZN(n585) );
  XNOR2_X1 U426 ( .A(n432), .B(KEYINPUT6), .ZN(n650) );
  NOR2_X1 U427 ( .A1(n434), .A2(n725), .ZN(n608) );
  XNOR2_X1 U428 ( .A(n715), .B(n483), .ZN(n434) );
  NAND2_X1 U429 ( .A1(n376), .A2(n647), .ZN(n491) );
  XNOR2_X1 U430 ( .A(n484), .B(n584), .ZN(n715) );
  NOR2_X1 U431 ( .A1(n673), .A2(G902), .ZN(n484) );
  XOR2_X1 U432 ( .A(n752), .B(KEYINPUT59), .Z(n754) );
  AND2_X1 U433 ( .A1(G224), .A2(n531), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n429), .B(KEYINPUT67), .ZN(n580) );
  INV_X1 U435 ( .A(n461), .ZN(n366) );
  NAND2_X1 U436 ( .A1(n779), .A2(n765), .ZN(n707) );
  NOR2_X1 U437 ( .A1(n600), .A2(n351), .ZN(n367) );
  NOR2_X1 U438 ( .A1(G953), .A2(G237), .ZN(n577) );
  XNOR2_X1 U439 ( .A(G125), .B(G146), .ZN(n545) );
  XNOR2_X1 U440 ( .A(n525), .B(n400), .ZN(n526) );
  XNOR2_X1 U441 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n524) );
  XNOR2_X1 U442 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n643) );
  INV_X1 U443 ( .A(KEYINPUT91), .ZN(n570) );
  INV_X1 U444 ( .A(G116), .ZN(n509) );
  INV_X1 U445 ( .A(KEYINPUT3), .ZN(n510) );
  XNOR2_X1 U446 ( .A(n555), .B(n556), .ZN(n426) );
  INV_X1 U447 ( .A(n752), .ZN(n391) );
  INV_X1 U448 ( .A(n705), .ZN(n508) );
  XNOR2_X1 U449 ( .A(n658), .B(n657), .ZN(n401) );
  OR2_X1 U450 ( .A1(n430), .A2(n476), .ZN(n493) );
  XNOR2_X1 U451 ( .A(n395), .B(n505), .ZN(n728) );
  INV_X1 U452 ( .A(KEYINPUT107), .ZN(n505) );
  NOR2_X1 U453 ( .A1(n724), .A2(n725), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n582), .B(n583), .ZN(n673) );
  XNOR2_X1 U455 ( .A(n587), .B(n368), .ZN(n582) );
  XNOR2_X1 U456 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U457 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U458 ( .A(n588), .B(G104), .ZN(n393) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(G143), .Z(n541) );
  XNOR2_X1 U460 ( .A(n431), .B(n776), .ZN(n668) );
  XNOR2_X1 U461 ( .A(n421), .B(n420), .ZN(n431) );
  XNOR2_X1 U462 ( .A(n589), .B(n590), .ZN(n420) );
  XNOR2_X1 U463 ( .A(n368), .B(n422), .ZN(n421) );
  NAND2_X1 U464 ( .A1(n499), .A2(n498), .ZN(n497) );
  NAND2_X1 U465 ( .A1(n503), .A2(n374), .ZN(n498) );
  NAND2_X1 U466 ( .A1(n502), .A2(n500), .ZN(n499) );
  XNOR2_X1 U467 ( .A(n523), .B(n522), .ZN(n771) );
  XNOR2_X1 U468 ( .A(n576), .B(n515), .ZN(n523) );
  XNOR2_X1 U469 ( .A(n526), .B(n398), .ZN(n453) );
  NAND2_X1 U470 ( .A1(n501), .A2(n399), .ZN(n398) );
  NAND2_X1 U471 ( .A1(n500), .A2(n374), .ZN(n399) );
  NAND2_X1 U472 ( .A1(n502), .A2(n503), .ZN(n501) );
  INV_X1 U473 ( .A(n725), .ZN(n470) );
  NAND2_X1 U474 ( .A1(n699), .A2(KEYINPUT40), .ZN(n447) );
  INV_X1 U475 ( .A(KEYINPUT36), .ZN(n467) );
  INV_X1 U476 ( .A(KEYINPUT1), .ZN(n594) );
  NAND2_X1 U477 ( .A1(n737), .A2(n418), .ZN(n417) );
  NOR2_X1 U478 ( .A1(n603), .A2(n434), .ZN(n606) );
  NAND2_X1 U479 ( .A1(n461), .A2(KEYINPUT2), .ZN(n460) );
  NAND2_X1 U480 ( .A1(n456), .A2(n455), .ZN(n454) );
  XNOR2_X1 U481 ( .A(n472), .B(n471), .ZN(n758) );
  XNOR2_X1 U482 ( .A(n538), .B(n534), .ZN(n471) );
  XNOR2_X1 U483 ( .A(n536), .B(n473), .ZN(n472) );
  NOR2_X1 U484 ( .A1(n695), .A2(n375), .ZN(n384) );
  NAND2_X1 U485 ( .A1(n371), .A2(n389), .ZN(n388) );
  NAND2_X1 U486 ( .A1(n386), .A2(n383), .ZN(n382) );
  NAND2_X1 U487 ( .A1(n388), .A2(n387), .ZN(n386) );
  AND2_X1 U488 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U489 ( .A(KEYINPUT47), .ZN(n387) );
  NAND2_X1 U490 ( .A1(n496), .A2(n494), .ZN(n476) );
  INV_X1 U491 ( .A(KEYINPUT82), .ZN(n494) );
  INV_X1 U492 ( .A(KEYINPUT4), .ZN(n429) );
  NAND2_X1 U493 ( .A1(n466), .A2(n426), .ZN(n713) );
  XNOR2_X1 U494 ( .A(n581), .B(n580), .ZN(n587) );
  XNOR2_X1 U495 ( .A(G110), .B(G119), .ZN(n558) );
  XNOR2_X1 U496 ( .A(G140), .B(G128), .ZN(n561) );
  XNOR2_X1 U497 ( .A(n537), .B(G134), .ZN(n581) );
  XNOR2_X1 U498 ( .A(n591), .B(KEYINPUT74), .ZN(n422) );
  INV_X1 U499 ( .A(G146), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n587), .B(n588), .ZN(n776) );
  XNOR2_X1 U501 ( .A(n521), .B(n520), .ZN(n589) );
  XNOR2_X1 U502 ( .A(G110), .B(G104), .ZN(n520) );
  NAND2_X1 U503 ( .A1(n512), .A2(n511), .ZN(n514) );
  INV_X1 U504 ( .A(n374), .ZN(n502) );
  INV_X1 U505 ( .A(n545), .ZN(n503) );
  INV_X1 U506 ( .A(n503), .ZN(n500) );
  NAND2_X1 U507 ( .A1(n728), .A2(n376), .ZN(n394) );
  AND2_X1 U508 ( .A1(n642), .A2(n643), .ZN(n418) );
  XNOR2_X1 U509 ( .A(n426), .B(n425), .ZN(n647) );
  INV_X1 U510 ( .A(KEYINPUT94), .ZN(n425) );
  XNOR2_X1 U511 ( .A(n475), .B(KEYINPUT72), .ZN(n404) );
  NOR2_X1 U512 ( .A1(n710), .A2(n709), .ZN(n475) );
  OR2_X1 U513 ( .A1(G902), .A2(G237), .ZN(n529) );
  NOR2_X1 U514 ( .A1(n610), .A2(n426), .ZN(n574) );
  XNOR2_X1 U515 ( .A(KEYINPUT13), .B(G475), .ZN(n488) );
  NAND2_X1 U516 ( .A1(n391), .A2(n390), .ZN(n489) );
  INV_X1 U517 ( .A(G902), .ZN(n390) );
  NAND2_X1 U518 ( .A1(n660), .A2(n647), .ZN(n709) );
  INV_X1 U519 ( .A(KEYINPUT81), .ZN(n506) );
  XNOR2_X1 U520 ( .A(n409), .B(KEYINPUT45), .ZN(n765) );
  NOR2_X1 U521 ( .A1(n492), .A2(n370), .ZN(n408) );
  XNOR2_X1 U522 ( .A(n535), .B(n533), .ZN(n473) );
  XOR2_X1 U523 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n535) );
  XNOR2_X1 U524 ( .A(n539), .B(n474), .ZN(n622) );
  XNOR2_X1 U525 ( .A(KEYINPUT98), .B(G478), .ZN(n474) );
  NOR2_X1 U526 ( .A1(G902), .A2(n758), .ZN(n539) );
  INV_X1 U527 ( .A(KEYINPUT100), .ZN(n483) );
  INV_X1 U528 ( .A(n660), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n675), .B(n674), .ZN(n677) );
  XNOR2_X1 U530 ( .A(n424), .B(n423), .ZN(n761) );
  XNOR2_X1 U531 ( .A(n564), .B(n566), .ZN(n424) );
  XNOR2_X1 U532 ( .A(n392), .B(n369), .ZN(n752) );
  XNOR2_X1 U533 ( .A(n372), .B(n393), .ZN(n392) );
  NAND2_X1 U534 ( .A1(n442), .A2(n441), .ZN(n439) );
  AND2_X1 U535 ( .A1(n444), .A2(n443), .ZN(n440) );
  NOR2_X1 U536 ( .A1(n436), .A2(n377), .ZN(n441) );
  NAND2_X1 U537 ( .A1(n446), .A2(n445), .ZN(n437) );
  NOR2_X1 U538 ( .A1(n699), .A2(KEYINPUT40), .ZN(n445) );
  XNOR2_X1 U539 ( .A(n599), .B(n467), .ZN(n600) );
  NAND2_X1 U540 ( .A1(n412), .A2(n411), .ZN(n410) );
  XNOR2_X1 U541 ( .A(n381), .B(KEYINPUT76), .ZN(n653) );
  OR2_X1 U542 ( .A1(n652), .A2(n660), .ZN(n381) );
  XNOR2_X1 U543 ( .A(n758), .B(n757), .ZN(n486) );
  INV_X1 U544 ( .A(n762), .ZN(n670) );
  XOR2_X1 U545 ( .A(n544), .B(n557), .Z(n369) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(n621) );
  AND2_X1 U547 ( .A1(n641), .A2(n640), .ZN(n370) );
  NAND2_X1 U548 ( .A1(n697), .A2(n640), .ZN(n371) );
  XOR2_X1 U549 ( .A(n541), .B(n540), .Z(n372) );
  XOR2_X1 U550 ( .A(G137), .B(G131), .Z(n373) );
  AND2_X1 U551 ( .A1(n727), .A2(KEYINPUT77), .ZN(n375) );
  AND2_X1 U552 ( .A1(n621), .A2(n622), .ZN(n376) );
  XNOR2_X1 U553 ( .A(G137), .B(KEYINPUT68), .ZN(n590) );
  XOR2_X1 U554 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n377) );
  XNOR2_X1 U555 ( .A(n394), .B(n602), .ZN(n722) );
  XOR2_X1 U556 ( .A(n668), .B(n667), .Z(n378) );
  NAND2_X1 U557 ( .A1(KEYINPUT44), .A2(KEYINPUT82), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n665), .A2(KEYINPUT79), .ZN(n379) );
  AND2_X1 U559 ( .A1(n666), .A2(n459), .ZN(n380) );
  INV_X1 U560 ( .A(n788), .ZN(n402) );
  XNOR2_X1 U561 ( .A(n655), .B(KEYINPUT32), .ZN(n788) );
  NAND2_X1 U562 ( .A1(n408), .A2(n405), .ZN(n409) );
  XNOR2_X1 U563 ( .A(n575), .B(n373), .ZN(n462) );
  INV_X1 U564 ( .A(n707), .ZN(n457) );
  NOR2_X1 U565 ( .A1(n631), .A2(n610), .ZN(n611) );
  XNOR2_X1 U566 ( .A(n573), .B(n572), .ZN(n712) );
  INV_X1 U567 ( .A(n777), .ZN(n423) );
  NAND2_X1 U568 ( .A1(n627), .A2(KEYINPUT47), .ZN(n385) );
  INV_X1 U569 ( .A(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U570 ( .A(n396), .B(n397), .ZN(n400) );
  INV_X1 U571 ( .A(n537), .ZN(n396) );
  XNOR2_X2 U572 ( .A(KEYINPUT66), .B(G101), .ZN(n397) );
  XNOR2_X2 U573 ( .A(G128), .B(G143), .ZN(n537) );
  INV_X1 U574 ( .A(n463), .ZN(n690) );
  NAND2_X1 U575 ( .A1(n495), .A2(n401), .ZN(n407) );
  NAND2_X1 U576 ( .A1(n609), .A2(n403), .ZN(n631) );
  NAND2_X1 U577 ( .A1(n607), .A2(n403), .ZN(n436) );
  NAND2_X1 U578 ( .A1(n404), .A2(n662), .ZN(n433) );
  NAND2_X1 U579 ( .A1(n404), .A2(n432), .ZN(n718) );
  NAND2_X1 U580 ( .A1(n468), .A2(KEYINPUT44), .ZN(n406) );
  INV_X1 U581 ( .A(n643), .ZN(n411) );
  INV_X1 U582 ( .A(n737), .ZN(n412) );
  NOR2_X1 U583 ( .A1(n416), .A2(n415), .ZN(n414) );
  INV_X1 U584 ( .A(n644), .ZN(n415) );
  NOR2_X1 U585 ( .A1(n642), .A2(n643), .ZN(n416) );
  XNOR2_X2 U586 ( .A(n419), .B(n645), .ZN(n430) );
  XNOR2_X1 U587 ( .A(n557), .B(n590), .ZN(n777) );
  NAND2_X1 U588 ( .A1(n665), .A2(G234), .ZN(n554) );
  XNOR2_X2 U589 ( .A(n427), .B(KEYINPUT86), .ZN(n665) );
  XNOR2_X2 U590 ( .A(G902), .B(KEYINPUT15), .ZN(n427) );
  NOR2_X1 U591 ( .A1(n436), .A2(n428), .ZN(n697) );
  XNOR2_X1 U592 ( .A(n618), .B(n617), .ZN(n428) );
  NAND2_X1 U593 ( .A1(n430), .A2(KEYINPUT82), .ZN(n656) );
  NOR2_X1 U594 ( .A1(n430), .A2(n477), .ZN(n495) );
  XNOR2_X1 U595 ( .A(n430), .B(n789), .ZN(G24) );
  BUF_X2 U596 ( .A(n715), .Z(n432) );
  XNOR2_X2 U597 ( .A(n433), .B(KEYINPUT33), .ZN(n737) );
  NAND2_X1 U598 ( .A1(n493), .A2(n664), .ZN(n492) );
  NAND2_X1 U599 ( .A1(n707), .A2(KEYINPUT79), .ZN(n458) );
  AND2_X1 U600 ( .A1(n434), .A2(n466), .ZN(n465) );
  NAND2_X1 U601 ( .A1(n436), .A2(n377), .ZN(n443) );
  NAND2_X1 U602 ( .A1(n504), .A2(n792), .ZN(n616) );
  INV_X1 U603 ( .A(n722), .ZN(n442) );
  NAND2_X1 U604 ( .A1(n722), .A2(n377), .ZN(n444) );
  INV_X1 U605 ( .A(n629), .ZN(n446) );
  NAND2_X1 U606 ( .A1(n629), .A2(KEYINPUT40), .ZN(n448) );
  NAND2_X1 U607 ( .A1(n450), .A2(n771), .ZN(n449) );
  XNOR2_X1 U608 ( .A(n526), .B(n497), .ZN(n450) );
  INV_X1 U609 ( .A(n771), .ZN(n452) );
  NAND2_X1 U610 ( .A1(n747), .A2(n665), .ZN(n528) );
  NAND2_X1 U611 ( .A1(n457), .A2(n379), .ZN(n455) );
  NAND2_X1 U612 ( .A1(n665), .A2(KEYINPUT79), .ZN(n459) );
  INV_X1 U613 ( .A(n707), .ZN(n461) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n630) );
  XNOR2_X1 U615 ( .A(n659), .B(n649), .ZN(n464) );
  XNOR2_X1 U616 ( .A(n576), .B(n462), .ZN(n579) );
  NOR2_X2 U617 ( .A1(n654), .A2(n651), .ZN(n659) );
  NAND2_X1 U618 ( .A1(n464), .A2(n465), .ZN(n463) );
  NAND2_X1 U619 ( .A1(n696), .A2(n470), .ZN(n469) );
  NAND2_X1 U620 ( .A1(n658), .A2(n656), .ZN(n468) );
  NAND2_X1 U621 ( .A1(n482), .A2(n628), .ZN(n481) );
  INV_X1 U622 ( .A(n496), .ZN(n477) );
  NAND2_X1 U623 ( .A1(n479), .A2(n508), .ZN(n507) );
  XNOR2_X1 U624 ( .A(n481), .B(n480), .ZN(n479) );
  INV_X1 U625 ( .A(KEYINPUT48), .ZN(n480) );
  NOR2_X1 U626 ( .A1(n485), .A2(n762), .ZN(G63) );
  XNOR2_X1 U627 ( .A(n487), .B(n486), .ZN(n485) );
  NAND2_X1 U628 ( .A1(n759), .A2(G478), .ZN(n487) );
  INV_X1 U629 ( .A(n696), .ZN(n699) );
  XNOR2_X1 U630 ( .A(n504), .B(G137), .ZN(G39) );
  NOR2_X1 U631 ( .A1(n625), .A2(n725), .ZN(n618) );
  INV_X1 U632 ( .A(KEYINPUT64), .ZN(n614) );
  INV_X1 U633 ( .A(KEYINPUT23), .ZN(n560) );
  XNOR2_X1 U634 ( .A(n608), .B(KEYINPUT30), .ZN(n612) );
  INV_X1 U635 ( .A(KEYINPUT22), .ZN(n648) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  INV_X1 U637 ( .A(KEYINPUT63), .ZN(n679) );
  NAND2_X1 U638 ( .A1(n509), .A2(KEYINPUT3), .ZN(n512) );
  NAND2_X1 U639 ( .A1(n510), .A2(G116), .ZN(n511) );
  XNOR2_X1 U640 ( .A(G122), .B(KEYINPUT16), .ZN(n515) );
  INV_X1 U641 ( .A(G107), .ZN(n516) );
  NAND2_X1 U642 ( .A1(n516), .A2(KEYINPUT87), .ZN(n519) );
  INV_X1 U643 ( .A(KEYINPUT87), .ZN(n517) );
  NAND2_X1 U644 ( .A1(n517), .A2(G107), .ZN(n518) );
  NAND2_X1 U645 ( .A1(n519), .A2(n518), .ZN(n521) );
  INV_X1 U646 ( .A(n589), .ZN(n522) );
  XNOR2_X1 U647 ( .A(n524), .B(n580), .ZN(n525) );
  NAND2_X1 U648 ( .A1(n529), .A2(G210), .ZN(n527) );
  XNOR2_X2 U649 ( .A(n528), .B(n527), .ZN(n625) );
  XOR2_X1 U650 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n596) );
  NAND2_X1 U651 ( .A1(G214), .A2(n529), .ZN(n530) );
  XOR2_X1 U652 ( .A(KEYINPUT88), .B(n530), .Z(n725) );
  NAND2_X1 U653 ( .A1(G234), .A2(n531), .ZN(n532) );
  XOR2_X1 U654 ( .A(KEYINPUT8), .B(n532), .Z(n565) );
  NAND2_X1 U655 ( .A1(G217), .A2(n565), .ZN(n536) );
  XOR2_X1 U656 ( .A(KEYINPUT9), .B(G116), .Z(n534) );
  XNOR2_X1 U657 ( .A(G122), .B(G107), .ZN(n533) );
  INV_X1 U658 ( .A(n581), .ZN(n538) );
  XOR2_X1 U659 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n543) );
  NAND2_X1 U660 ( .A1(n577), .A2(G214), .ZN(n542) );
  XNOR2_X1 U661 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U662 ( .A(G140), .B(G131), .Z(n588) );
  XNOR2_X1 U663 ( .A(KEYINPUT10), .B(n545), .ZN(n557) );
  INV_X1 U664 ( .A(n621), .ZN(n619) );
  NAND2_X1 U665 ( .A1(n622), .A2(n619), .ZN(n546) );
  XNOR2_X1 U666 ( .A(n546), .B(KEYINPUT99), .ZN(n696) );
  NAND2_X1 U667 ( .A1(G237), .A2(G234), .ZN(n547) );
  XNOR2_X1 U668 ( .A(n547), .B(KEYINPUT14), .ZN(n549) );
  NAND2_X1 U669 ( .A1(n549), .A2(G952), .ZN(n548) );
  XOR2_X1 U670 ( .A(KEYINPUT89), .B(n548), .Z(n736) );
  NOR2_X1 U671 ( .A1(G953), .A2(n736), .ZN(n634) );
  NAND2_X1 U672 ( .A1(G902), .A2(n549), .ZN(n550) );
  XOR2_X1 U673 ( .A(KEYINPUT90), .B(n550), .Z(n551) );
  NAND2_X1 U674 ( .A1(G953), .A2(n551), .ZN(n632) );
  NOR2_X1 U675 ( .A1(G900), .A2(n632), .ZN(n552) );
  XNOR2_X1 U676 ( .A(n552), .B(KEYINPUT102), .ZN(n553) );
  NOR2_X1 U677 ( .A1(n634), .A2(n553), .ZN(n610) );
  XOR2_X1 U678 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n556) );
  XNOR2_X1 U679 ( .A(n554), .B(KEYINPUT20), .ZN(n567) );
  NAND2_X1 U680 ( .A1(n567), .A2(G221), .ZN(n555) );
  XOR2_X1 U681 ( .A(KEYINPUT24), .B(KEYINPUT73), .Z(n559) );
  XNOR2_X1 U682 ( .A(n559), .B(n558), .ZN(n563) );
  NAND2_X1 U683 ( .A1(G221), .A2(n565), .ZN(n566) );
  NOR2_X1 U684 ( .A1(n761), .A2(G902), .ZN(n573) );
  XOR2_X1 U685 ( .A(KEYINPUT92), .B(KEYINPUT25), .Z(n569) );
  NAND2_X1 U686 ( .A1(n567), .A2(G217), .ZN(n568) );
  XNOR2_X1 U687 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U688 ( .A1(n574), .A2(n712), .ZN(n603) );
  XOR2_X1 U689 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n575) );
  NAND2_X1 U690 ( .A1(n577), .A2(G210), .ZN(n578) );
  XNOR2_X1 U691 ( .A(n579), .B(n578), .ZN(n583) );
  NAND2_X1 U692 ( .A1(G227), .A2(n531), .ZN(n591) );
  XNOR2_X1 U693 ( .A(KEYINPUT69), .B(G469), .ZN(n592) );
  NAND2_X1 U694 ( .A1(n598), .A2(n351), .ZN(n595) );
  XNOR2_X1 U695 ( .A(n596), .B(n595), .ZN(n597) );
  NOR2_X1 U696 ( .A1(n601), .A2(n597), .ZN(n705) );
  XOR2_X1 U697 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n602) );
  XOR2_X1 U698 ( .A(KEYINPUT105), .B(KEYINPUT28), .Z(n604) );
  XNOR2_X1 U699 ( .A(KEYINPUT106), .B(n604), .ZN(n605) );
  XNOR2_X1 U700 ( .A(n606), .B(n605), .ZN(n607) );
  INV_X1 U701 ( .A(n709), .ZN(n609) );
  NAND2_X1 U702 ( .A1(n612), .A2(n611), .ZN(n620) );
  XNOR2_X1 U703 ( .A(KEYINPUT70), .B(KEYINPUT39), .ZN(n613) );
  XNOR2_X1 U704 ( .A(n616), .B(n615), .ZN(n628) );
  XOR2_X1 U705 ( .A(KEYINPUT65), .B(KEYINPUT19), .Z(n617) );
  NOR2_X1 U706 ( .A1(n619), .A2(n622), .ZN(n691) );
  INV_X1 U707 ( .A(n691), .ZN(n702) );
  NAND2_X1 U708 ( .A1(n702), .A2(n699), .ZN(n727) );
  XNOR2_X1 U709 ( .A(n727), .B(KEYINPUT78), .ZN(n640) );
  INV_X1 U710 ( .A(n620), .ZN(n623) );
  NOR2_X1 U711 ( .A1(n622), .A2(n621), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n623), .A2(n644), .ZN(n624) );
  NOR2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n695) );
  OR2_X1 U714 ( .A1(KEYINPUT77), .A2(n727), .ZN(n626) );
  NAND2_X1 U715 ( .A1(n626), .A2(n697), .ZN(n627) );
  NOR2_X1 U716 ( .A1(n629), .A2(n702), .ZN(n704) );
  NOR2_X2 U717 ( .A1(n630), .A2(n704), .ZN(n779) );
  NOR2_X1 U718 ( .A1(n432), .A2(n631), .ZN(n638) );
  NOR2_X1 U719 ( .A1(G898), .A2(n632), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n635) );
  INV_X1 U721 ( .A(KEYINPUT0), .ZN(n636) );
  INV_X1 U722 ( .A(n646), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n638), .A2(n642), .ZN(n684) );
  NOR2_X1 U724 ( .A1(n718), .A2(n646), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(KEYINPUT31), .ZN(n701) );
  NAND2_X1 U726 ( .A1(n684), .A2(n701), .ZN(n641) );
  INV_X1 U727 ( .A(n650), .ZN(n662) );
  XNOR2_X1 U728 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n645) );
  INV_X1 U729 ( .A(KEYINPUT101), .ZN(n649) );
  INV_X1 U730 ( .A(n710), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  INV_X1 U733 ( .A(KEYINPUT83), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n681) );
  NOR2_X1 U736 ( .A1(KEYINPUT44), .A2(KEYINPUT82), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n681), .A2(n663), .ZN(n664) );
  INV_X1 U738 ( .A(KEYINPUT2), .ZN(n708) );
  OR2_X1 U739 ( .A1(n708), .A2(n665), .ZN(n666) );
  NAND2_X1 U740 ( .A1(n759), .A2(G469), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n667) );
  XNOR2_X1 U742 ( .A(n669), .B(n378), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT119), .ZN(G54) );
  XNOR2_X1 U745 ( .A(KEYINPUT85), .B(KEYINPUT111), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n350), .B(KEYINPUT62), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n759), .A2(G472), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(G57) );
  XOR2_X1 U749 ( .A(G101), .B(n681), .Z(n682) );
  XNOR2_X1 U750 ( .A(KEYINPUT112), .B(n682), .ZN(G3) );
  NOR2_X1 U751 ( .A1(n699), .A2(n684), .ZN(n683) );
  XOR2_X1 U752 ( .A(G104), .B(n683), .Z(G6) );
  NOR2_X1 U753 ( .A1(n702), .A2(n684), .ZN(n689) );
  XOR2_X1 U754 ( .A(KEYINPUT114), .B(KEYINPUT27), .Z(n686) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT26), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U757 ( .A(KEYINPUT113), .B(n687), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n689), .B(n688), .ZN(G9) );
  XOR2_X1 U759 ( .A(n690), .B(G110), .Z(G12) );
  XOR2_X1 U760 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n693) );
  NAND2_X1 U761 ( .A1(n697), .A2(n691), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U763 ( .A(G128), .B(n694), .Z(G30) );
  XOR2_X1 U764 ( .A(G143), .B(n695), .Z(G45) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n698), .B(G146), .ZN(G48) );
  NOR2_X1 U767 ( .A1(n699), .A2(n701), .ZN(n700) );
  XOR2_X1 U768 ( .A(G113), .B(n700), .Z(G15) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U770 ( .A(G116), .B(n703), .Z(G18) );
  XOR2_X1 U771 ( .A(G134), .B(n704), .Z(G36) );
  XOR2_X1 U772 ( .A(G140), .B(n705), .Z(n706) );
  XNOR2_X1 U773 ( .A(KEYINPUT116), .B(n706), .ZN(G42) );
  XNOR2_X1 U774 ( .A(n708), .B(n366), .ZN(n741) );
  NAND2_X1 U775 ( .A1(n351), .A2(n709), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT50), .ZN(n717) );
  XNOR2_X1 U777 ( .A(KEYINPUT49), .B(n713), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n432), .A2(n714), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U781 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n720) );
  XNOR2_X1 U782 ( .A(n721), .B(n720), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n723), .A2(n442), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U785 ( .A1(n726), .A2(n376), .ZN(n730) );
  NAND2_X1 U786 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n352), .A2(n731), .ZN(n732) );
  NAND2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U790 ( .A(KEYINPUT52), .B(n734), .Z(n735) );
  NOR2_X1 U791 ( .A1(n736), .A2(n735), .ZN(n739) );
  AND2_X1 U792 ( .A1(n352), .A2(n442), .ZN(n738) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U795 ( .A1(n742), .A2(G953), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n743), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U797 ( .A(KEYINPUT55), .B(KEYINPUT84), .Z(n745) );
  XNOR2_X1 U798 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n745), .B(n744), .ZN(n746) );
  XOR2_X1 U800 ( .A(n747), .B(n746), .Z(n749) );
  NAND2_X1 U801 ( .A1(n759), .A2(G210), .ZN(n748) );
  XNOR2_X1 U802 ( .A(n751), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U803 ( .A1(n759), .A2(G475), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n756), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U805 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n757) );
  XNOR2_X1 U806 ( .A(n760), .B(n761), .ZN(n763) );
  XNOR2_X1 U807 ( .A(n764), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U808 ( .A1(n531), .A2(n765), .ZN(n770) );
  NAND2_X1 U809 ( .A1(G953), .A2(G224), .ZN(n766) );
  XNOR2_X1 U810 ( .A(KEYINPUT61), .B(n766), .ZN(n767) );
  NAND2_X1 U811 ( .A1(n767), .A2(G898), .ZN(n768) );
  XOR2_X1 U812 ( .A(KEYINPUT123), .B(n768), .Z(n769) );
  NAND2_X1 U813 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U814 ( .A(n771), .B(G101), .ZN(n773) );
  NOR2_X1 U815 ( .A1(n531), .A2(G898), .ZN(n772) );
  NOR2_X1 U816 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U817 ( .A(n775), .B(n774), .ZN(G69) );
  XNOR2_X1 U818 ( .A(n776), .B(n777), .ZN(n778) );
  XNOR2_X1 U819 ( .A(n778), .B(KEYINPUT124), .ZN(n782) );
  XNOR2_X1 U820 ( .A(n782), .B(n779), .ZN(n780) );
  NOR2_X1 U821 ( .A1(G953), .A2(n780), .ZN(n781) );
  XNOR2_X1 U822 ( .A(KEYINPUT125), .B(n781), .ZN(n786) );
  XNOR2_X1 U823 ( .A(G227), .B(n782), .ZN(n783) );
  NAND2_X1 U824 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U825 ( .A1(n784), .A2(G953), .ZN(n785) );
  NAND2_X1 U826 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U827 ( .A(n787), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U828 ( .A(G119), .B(n788), .Z(G21) );
  XNOR2_X1 U829 ( .A(G122), .B(KEYINPUT127), .ZN(n789) );
  XNOR2_X1 U830 ( .A(G125), .B(KEYINPUT37), .ZN(n791) );
  XNOR2_X1 U831 ( .A(n791), .B(n790), .ZN(G27) );
  XNOR2_X1 U832 ( .A(n792), .B(G131), .ZN(G33) );
endmodule

