//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G58), .A2(G232), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G77), .A2(G244), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G50), .A2(G226), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n210), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n216), .B1(new_n215), .B2(new_n214), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(G257), .A2(G264), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n224), .A2(new_n208), .A3(new_n225), .ZN(new_n226));
  AND3_X1   g0026(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n227));
  AOI21_X1  g0027(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI22_X1  g0034(.A1(new_n226), .A2(KEYINPUT0), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n222), .B(new_n235), .C1(KEYINPUT0), .C2(new_n226), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT7), .B1(new_n257), .B2(new_n230), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G159), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n230), .A2(new_n260), .A3(KEYINPUT69), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT69), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G20), .B2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G58), .A2(G68), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n230), .B1(new_n232), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n265), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n220), .B2(new_n260), .ZN(new_n279));
  NAND4_X1  g0079(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n229), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n261), .A2(new_n230), .A3(new_n262), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n263), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n273), .B1(new_n286), .B2(G68), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(KEYINPUT16), .A3(new_n271), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n277), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(G223), .B2(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G226), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(new_n260), .B2(new_n207), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n229), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n293), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G1), .A2(G13), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n299), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(new_n291), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G232), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(G190), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n301), .ZN(new_n309));
  INV_X1    g0109(.A(new_n293), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G200), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n290), .A2(G20), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n281), .A2(new_n229), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G1), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n315), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT80), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n317), .A2(KEYINPUT80), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n289), .A2(new_n308), .A3(new_n312), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT17), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  AOI21_X1  g0130(.A(G169), .B1(new_n302), .B2(new_n307), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n289), .B2(new_n326), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n302), .A2(new_n333), .A3(new_n307), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n332), .A2(KEYINPUT18), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT18), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n329), .B(new_n330), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n294), .A2(G232), .A3(G1698), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n294), .A2(G226), .A3(new_n296), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n260), .C2(new_n217), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n293), .B1(new_n341), .B2(new_n301), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n306), .A2(G238), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n342), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT14), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n341), .A2(new_n301), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(new_n310), .A3(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G179), .A3(new_n346), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n343), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n346), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G169), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n350), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G68), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(G77), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n230), .A2(G33), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n267), .A2(new_n269), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n361), .B1(new_n362), .B2(new_n363), .C1(new_n364), .C2(new_n202), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n282), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT11), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n314), .A2(new_n360), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n319), .A2(G20), .A3(new_n360), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n359), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n353), .A2(G190), .A3(new_n346), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT79), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT79), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n353), .A2(new_n377), .A3(G190), .A4(new_n346), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n373), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G200), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n355), .B2(new_n346), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G20), .A2(G77), .ZN(new_n384));
  OR2_X1    g0184(.A1(KEYINPUT15), .A2(G87), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT15), .A2(G87), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT73), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(KEYINPUT73), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n384), .B1(new_n364), .B2(new_n315), .C1(new_n391), .C2(new_n363), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n314), .A2(KEYINPUT75), .A3(new_n362), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT75), .B1(new_n314), .B2(new_n362), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n282), .A2(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n320), .A2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT74), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n294), .A2(G232), .A3(new_n296), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n257), .A2(G107), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n294), .A2(KEYINPUT72), .A3(G232), .A4(new_n296), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n293), .B1(new_n405), .B2(new_n301), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n306), .A2(G244), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n333), .A3(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n398), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n338), .A2(new_n374), .A3(new_n383), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n203), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(G150), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n414), .B1(new_n315), .B2(new_n363), .C1(new_n364), .C2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n320), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n416), .A2(new_n282), .B1(new_n202), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n313), .A2(G50), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT70), .ZN(new_n420));
  INV_X1    g0220(.A(new_n282), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n320), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n296), .A2(G222), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G223), .A2(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n294), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n301), .B(new_n426), .C1(G77), .C2(new_n294), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n306), .A2(G226), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n310), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n423), .B1(new_n430), .B2(G169), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT71), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G179), .B2(new_n429), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n395), .B(new_n397), .C1(new_n408), .C2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n380), .B1(new_n406), .B2(new_n407), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT10), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n429), .A2(new_n434), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n418), .A2(new_n441), .A3(new_n422), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n418), .B2(new_n422), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n430), .A2(new_n380), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n444), .B2(KEYINPUT77), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n442), .B2(new_n443), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n438), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n442), .A2(new_n443), .A3(new_n449), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n451), .A2(new_n452), .A3(new_n439), .A4(new_n446), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n433), .B(new_n437), .C1(new_n448), .C2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(G238), .B(new_n296), .C1(new_n255), .C2(new_n256), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  OAI21_X1  g0256(.A(G244), .B1(new_n255), .B2(new_n256), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(new_n456), .C1(new_n457), .C2(new_n296), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n301), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n305), .B(G250), .C1(G1), .C2(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n460), .A2(new_n292), .A3(G1), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n459), .A2(G190), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n294), .A2(new_n230), .A3(G68), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n230), .B1(new_n260), .B2(new_n217), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n207), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT19), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT19), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n363), .B2(new_n217), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n465), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n282), .B1(new_n391), .B2(new_n417), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n290), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n281), .A2(new_n229), .A3(new_n320), .A4(new_n474), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n475), .A2(new_n207), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n464), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n462), .B1(new_n458), .B2(new_n301), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n380), .B1(new_n478), .B2(new_n461), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n319), .A2(G20), .A3(new_n481), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT25), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n230), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n294), .A2(new_n489), .A3(new_n230), .A4(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n230), .A2(G33), .A3(G116), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT23), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n493), .A2(new_n230), .A3(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT23), .B1(new_n481), .B2(G20), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n488), .B2(new_n490), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT24), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(new_n492), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n486), .B1(new_n503), .B2(new_n282), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n208), .A2(new_n296), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n218), .A2(G1698), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n255), .C2(new_n256), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G294), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n301), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT5), .B(G41), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n462), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n462), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n460), .A2(G1), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n514), .A2(new_n520), .B1(new_n304), .B2(new_n299), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G264), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n380), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n513), .A2(new_n434), .A3(new_n519), .A4(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n480), .B1(new_n504), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT85), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G179), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n391), .A2(KEYINPUT86), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n389), .A2(new_n532), .A3(new_n390), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n473), .B1(new_n534), .B2(new_n475), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n409), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n333), .A4(new_n461), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n530), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n409), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n513), .A2(new_n333), .A3(new_n519), .A4(new_n522), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n421), .B1(new_n499), .B2(new_n502), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n486), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n527), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G264), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n294), .B(new_n545), .C1(new_n218), .C2(G1698), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n257), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n301), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT87), .B1(new_n521), .B2(G270), .ZN(new_n550));
  AND2_X1   g0350(.A1(KEYINPUT5), .A2(G41), .ZN(new_n551));
  NOR2_X1   g0351(.A1(KEYINPUT5), .A2(G41), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n520), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND4_X1   g0353(.A1(KEYINPUT87), .A2(new_n553), .A3(new_n305), .A4(G270), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n549), .B(new_n519), .C1(new_n550), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G20), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(G33), .B2(G283), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n260), .A2(G97), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n282), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n281), .A2(new_n229), .B1(new_n560), .B2(new_n559), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n558), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n475), .A2(G116), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n417), .A2(G116), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n564), .A2(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n544), .B1(new_n556), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n569), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n565), .A2(KEYINPUT20), .A3(new_n558), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT20), .B1(new_n565), .B2(new_n558), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n555), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n555), .A2(new_n333), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n575), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n571), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n555), .A2(new_n434), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G200), .B2(new_n555), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n581), .B2(new_n570), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n457), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n294), .A2(G250), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n296), .B1(new_n589), .B2(KEYINPUT4), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n583), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT4), .B1(new_n257), .B2(new_n208), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G1698), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n457), .A2(new_n585), .B1(G33), .B2(G283), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(KEYINPUT82), .A3(new_n594), .A4(new_n584), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n301), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n516), .A2(new_n518), .B1(new_n521), .B2(G257), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n481), .B1(new_n285), .B2(new_n263), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n217), .A2(new_n481), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n467), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n481), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n230), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n364), .A2(new_n362), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n600), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n421), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n475), .A2(G97), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n320), .A2(new_n217), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT81), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n610), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n596), .A2(new_n597), .A3(G190), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n599), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n598), .A2(new_n409), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n596), .A2(new_n597), .A3(new_n333), .ZN(new_n618));
  INV_X1    g0418(.A(new_n613), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n619), .A2(new_n611), .B1(new_n421), .B2(new_n607), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n616), .B2(new_n621), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n543), .B(new_n582), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n413), .A2(new_n454), .A3(new_n625), .ZN(G372));
  NOR2_X1   g0426(.A1(new_n413), .A2(new_n454), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n535), .B(new_n536), .C1(G179), .C2(new_n529), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n473), .A2(new_n476), .ZN(new_n629));
  INV_X1    g0429(.A(new_n529), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n464), .C1(new_n380), .C2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n538), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT26), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n527), .A2(new_n616), .A3(new_n621), .ZN(new_n634));
  INV_X1    g0434(.A(new_n542), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n579), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n628), .B(new_n633), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n631), .A2(new_n628), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n621), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n627), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n433), .ZN(new_n642));
  INV_X1    g0442(.A(new_n331), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT16), .B1(new_n287), .B2(new_n271), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n360), .B1(new_n285), .B2(new_n263), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n645), .A2(new_n276), .A3(new_n270), .A4(new_n273), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n644), .A2(new_n646), .A3(new_n421), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n324), .A2(new_n325), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n643), .B(new_n334), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n332), .A2(KEYINPUT18), .A3(new_n334), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n412), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n383), .A2(new_n654), .B1(new_n373), .B2(new_n359), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n330), .A2(new_n329), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n448), .A2(new_n453), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n642), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n641), .A2(new_n659), .ZN(G369));
  XOR2_X1   g0460(.A(KEYINPUT89), .B(KEYINPUT27), .Z(new_n661));
  NOR3_X1   g0461(.A1(new_n318), .A2(G1), .A3(G20), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n570), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n579), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n571), .A2(new_n576), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n581), .A2(new_n570), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(new_n578), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n673), .B2(new_n669), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n504), .A2(new_n526), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n667), .B1(new_n541), .B2(new_n486), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n501), .A2(new_n491), .A3(new_n492), .A4(new_n497), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n501), .B1(new_n500), .B2(new_n492), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n282), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(new_n485), .B1(new_n409), .B2(new_n523), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n675), .A2(new_n676), .B1(new_n680), .B2(new_n540), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n542), .A2(new_n667), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n674), .A2(G330), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n542), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n579), .A2(new_n668), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(G399));
  NOR2_X1   g0489(.A1(new_n224), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n468), .A2(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n233), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n616), .A2(new_n621), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT84), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n543), .A3(new_n582), .A4(new_n668), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n577), .A2(new_n522), .A3(new_n513), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n596), .A2(new_n630), .A3(new_n597), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n598), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n513), .A2(new_n522), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n707), .A2(new_n555), .A3(new_n333), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT30), .A4(new_n630), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT90), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n529), .B(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n523), .A2(new_n333), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n598), .A4(new_n555), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n705), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n714), .B2(new_n667), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n696), .B1(new_n701), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT26), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n621), .B2(new_n632), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n621), .A2(new_n638), .A3(new_n719), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT91), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n723), .B(new_n719), .C1(new_n621), .C2(new_n632), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n527), .A2(new_n616), .A3(new_n621), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n635), .B2(new_n579), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n671), .A2(KEYINPUT92), .A3(new_n542), .A4(new_n578), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n628), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT29), .B(new_n668), .C1(new_n725), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n668), .B1(new_n637), .B2(new_n639), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n718), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n695), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n318), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n691), .A2(G1), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n674), .B2(G330), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n674), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n224), .A2(new_n294), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n234), .A2(new_n460), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n744), .B(new_n745), .C1(new_n253), .C2(new_n460), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n294), .A2(G355), .A3(new_n223), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n747), .C1(G116), .C2(new_n223), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n229), .B1(G20), .B2(new_n409), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n740), .B(KEYINPUT93), .Z(new_n755));
  NOR2_X1   g0555(.A1(new_n230), .A2(new_n434), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n333), .A2(new_n380), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n380), .A2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n230), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G329), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n763), .A2(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n333), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n762), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n760), .B(new_n768), .C1(G311), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n756), .A2(new_n769), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G322), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n230), .B1(new_n765), .B2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G294), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n756), .A2(new_n761), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n257), .B1(new_n779), .B2(new_n547), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n757), .A2(new_n762), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n772), .A2(new_n775), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n758), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G50), .A2(new_n786), .B1(new_n771), .B2(G77), .ZN(new_n787));
  INV_X1    g0587(.A(new_n779), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G87), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n763), .A2(new_n481), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n787), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n781), .A2(new_n360), .B1(new_n776), .B2(new_n217), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT94), .ZN(new_n794));
  INV_X1    g0594(.A(new_n766), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n257), .B1(new_n796), .B2(KEYINPUT32), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n792), .A2(new_n794), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G58), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n773), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n785), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n755), .B1(new_n802), .B2(new_n749), .ZN(new_n803));
  INV_X1    g0603(.A(new_n752), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n754), .B(new_n803), .C1(new_n674), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n743), .A2(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n412), .A2(new_n667), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n398), .A2(new_n667), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n435), .B2(new_n436), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n412), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n733), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n668), .B(new_n810), .C1(new_n637), .C2(new_n639), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n718), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n718), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n814), .A2(new_n815), .A3(new_n741), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n763), .A2(new_n207), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n294), .B(new_n817), .C1(G283), .C2(new_n782), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n788), .A2(G107), .ZN(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n773), .A2(new_n820), .B1(new_n766), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G303), .B2(new_n786), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G116), .A2(new_n771), .B1(new_n777), .B2(G97), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n818), .A2(new_n819), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G143), .A2(new_n774), .B1(new_n782), .B2(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n827), .B2(new_n758), .C1(new_n266), .C2(new_n770), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT95), .Z(new_n829));
  OR2_X1    g0629(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n257), .B1(new_n795), .B2(G132), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  INV_X1    g0635(.A(new_n763), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G68), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n800), .B2(new_n776), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n779), .A2(new_n202), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n825), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n755), .B1(new_n842), .B2(new_n749), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n749), .A2(new_n750), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(G77), .B2(new_n845), .C1(new_n751), .C2(new_n810), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n816), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NAND2_X1  g0649(.A1(new_n289), .A2(new_n326), .ZN(new_n850));
  INV_X1    g0650(.A(new_n665), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n335), .A2(new_n336), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n656), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n332), .A2(new_n334), .B1(new_n850), .B2(new_n851), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT37), .B1(new_n856), .B2(new_n327), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n649), .A2(new_n852), .A3(new_n327), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n855), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n861), .B1(new_n337), .B2(new_n853), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n373), .B(new_n381), .C1(new_n376), .C2(new_n378), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n373), .B(new_n667), .C1(new_n869), .C2(new_n359), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n373), .A2(new_n667), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n374), .A2(new_n383), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n807), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n813), .A2(KEYINPUT98), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT98), .B1(new_n813), .B2(new_n874), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n868), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n374), .A2(new_n667), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT99), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n649), .A2(new_n852), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT100), .B1(new_n856), .B2(new_n327), .ZN(new_n884));
  AND4_X1   g0684(.A1(KEYINPUT100), .A2(new_n649), .A3(new_n327), .A4(new_n852), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n860), .B1(new_n856), .B2(new_n881), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT100), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n859), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n856), .A2(KEYINPUT100), .A3(new_n327), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n886), .A2(new_n855), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n864), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n867), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n866), .B2(new_n858), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n327), .B(KEYINPUT17), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n852), .B1(new_n653), .B2(new_n897), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n898), .A2(new_n864), .A3(new_n857), .A4(new_n861), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT39), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n880), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n653), .A2(new_n851), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n878), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n732), .A2(new_n627), .A3(new_n735), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n659), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(KEYINPUT102), .A2(KEYINPUT31), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n714), .A2(new_n667), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n714), .B2(new_n667), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n625), .A2(new_n667), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n811), .B1(new_n870), .B2(new_n872), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n910), .B(new_n911), .C1(new_n896), .C2(new_n899), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n911), .A2(new_n910), .A3(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n893), .A2(new_n867), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n627), .A2(new_n910), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n906), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n290), .B2(new_n738), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n272), .A2(G77), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n233), .A2(new_n922), .B1(G50), .B2(new_n360), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n318), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n603), .A2(new_n604), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n557), .B1(new_n925), .B2(KEYINPUT35), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n231), .C1(KEYINPUT35), .C2(new_n925), .ZN(new_n927));
  XOR2_X1   g0727(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n928));
  XNOR2_X1  g0728(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n924), .A3(new_n929), .ZN(G367));
  AOI22_X1  g0730(.A1(G58), .A2(new_n788), .B1(new_n774), .B2(G150), .ZN(new_n931));
  INV_X1    g0731(.A(G143), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n931), .B1(new_n827), .B2(new_n766), .C1(new_n932), .C2(new_n758), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n257), .B(new_n933), .C1(G77), .C2(new_n836), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n781), .A2(new_n266), .B1(new_n770), .B2(new_n202), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT110), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n934), .B(new_n936), .C1(new_n360), .C2(new_n776), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G303), .A2(new_n774), .B1(new_n771), .B2(G283), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n938), .B1(new_n821), .B2(new_n758), .C1(new_n939), .C2(new_n766), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G107), .B2(new_n777), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n836), .A2(G97), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n779), .B2(new_n557), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(new_n820), .C2(new_n781), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT109), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n942), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n294), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n755), .B1(new_n950), .B2(new_n749), .ZN(new_n951));
  INV_X1    g0751(.A(new_n744), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n753), .B1(new_n223), .B2(new_n391), .C1(new_n244), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n628), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n629), .A2(new_n668), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n638), .B2(new_n955), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n951), .B(new_n953), .C1(new_n804), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n739), .A2(G1), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n620), .A2(new_n667), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n616), .A2(new_n621), .A3(new_n962), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n617), .A2(new_n618), .A3(new_n620), .A4(new_n667), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n688), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n963), .A2(new_n964), .ZN(new_n969));
  INV_X1    g0769(.A(new_n682), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n579), .A2(new_n668), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n681), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n968), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n688), .A2(new_n965), .A3(new_n967), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n972), .A3(new_n960), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n966), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n684), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n683), .B(new_n971), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT108), .B1(new_n674), .B2(G330), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n684), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n976), .A2(KEYINPUT107), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n736), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n736), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n690), .B(KEYINPUT41), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n959), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n683), .A2(new_n965), .A3(new_n687), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT42), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n683), .A2(new_n965), .A3(KEYINPUT42), .A4(new_n687), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n621), .B1(new_n963), .B2(new_n542), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n990), .A2(new_n991), .B1(new_n668), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT103), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n957), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n993), .A2(KEYINPUT104), .A3(new_n997), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT104), .B1(new_n993), .B2(new_n997), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n684), .A2(new_n969), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n958), .B1(new_n987), .B2(new_n1008), .ZN(G387));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n777), .A2(G283), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n758), .A2(new_n1012), .B1(new_n781), .B2(new_n821), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT113), .Z(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n547), .B2(new_n770), .C1(new_n939), .C2(new_n773), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1011), .B1(new_n820), .B2(new_n779), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1010), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n294), .B1(new_n836), .B2(G116), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n766), .A2(new_n759), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1018), .A2(new_n1010), .A3(new_n1019), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G159), .A2(new_n786), .B1(new_n771), .B2(G68), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n315), .B2(new_n781), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n788), .A2(G77), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n795), .A2(G150), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n942), .A3(new_n1029), .A4(new_n294), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1027), .B1(KEYINPUT112), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n531), .A2(new_n533), .A3(new_n777), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(KEYINPUT112), .C2(new_n1030), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G50), .B2(new_n774), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n749), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n683), .A2(new_n804), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n315), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT111), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n692), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n360), .A2(new_n362), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(G45), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n744), .B1(new_n241), .B2(new_n460), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1043), .A2(new_n1044), .B1(G107), .B2(new_n223), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n692), .A2(new_n224), .A3(new_n257), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n755), .B(new_n1036), .C1(new_n753), .C2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1035), .A2(new_n1048), .B1(new_n959), .B2(new_n981), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n736), .A2(new_n981), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n690), .B1(new_n736), .B2(new_n981), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  XNOR2_X1  g0852(.A(new_n976), .B(new_n684), .ZN(new_n1053));
  OAI21_X1  g0853(.A(KEYINPUT115), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n736), .A2(new_n981), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n976), .B(new_n982), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT115), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n690), .A3(new_n984), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n969), .A2(new_n752), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n753), .B1(new_n217), .B2(new_n223), .C1(new_n250), .C2(new_n952), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n781), .A2(new_n547), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n770), .A2(new_n820), .B1(new_n766), .B2(new_n1012), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G283), .C2(new_n788), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n758), .A2(new_n939), .B1(new_n773), .B2(new_n821), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n294), .B1(new_n777), .B2(G116), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n791), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n782), .A2(G50), .B1(new_n771), .B2(new_n316), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n360), .B2(new_n779), .C1(new_n932), .C2(new_n766), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G77), .B2(new_n777), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n758), .A2(new_n415), .B1(new_n773), .B2(new_n266), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n294), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1074), .B2(new_n817), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n755), .B1(new_n1075), .B2(new_n749), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1060), .A2(new_n1061), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1053), .B2(new_n959), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1059), .A2(new_n1078), .ZN(G390));
  INV_X1    g0879(.A(KEYINPUT116), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n627), .A2(G330), .A3(new_n910), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n904), .A2(new_n1081), .A3(new_n659), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n876), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n813), .A2(KEYINPUT98), .A3(new_n874), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n810), .A2(G330), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n910), .A2(new_n873), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n701), .B2(new_n717), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n873), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n809), .A2(new_n412), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n668), .B(new_n1092), .C1(new_n725), .C2(new_n731), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n874), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n910), .A2(new_n1087), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n873), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1089), .A2(new_n873), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1080), .B(new_n1082), .C1(new_n1091), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1091), .A2(new_n1099), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1082), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT116), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n895), .A2(new_n900), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n880), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n915), .A2(new_n880), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1093), .A2(new_n874), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n873), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1088), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n880), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1105), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1098), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n880), .B(new_n915), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT117), .B1(new_n1104), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n691), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1123), .A2(new_n1094), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1080), .B1(new_n1124), .B2(new_n1082), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1101), .A2(KEYINPUT116), .A3(new_n1102), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n1111), .A4(new_n1117), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1119), .A2(new_n1122), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1113), .A2(new_n750), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n774), .A2(G116), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n789), .A2(new_n1132), .A3(new_n837), .A4(new_n257), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G107), .A2(new_n782), .B1(new_n795), .B2(G294), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n217), .B2(new_n770), .C1(new_n764), .C2(new_n758), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(G77), .C2(new_n777), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n779), .A2(new_n415), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n266), .B2(new_n776), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n770), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n795), .A2(G125), .ZN(new_n1143));
  INV_X1    g0943(.A(G132), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n773), .C1(new_n827), .C2(new_n781), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n294), .B1(new_n763), .B2(new_n202), .C1(new_n1146), .C2(new_n758), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1140), .A2(new_n1142), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n749), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n755), .B1(new_n315), .B2(new_n844), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT118), .Z(new_n1151));
  AND3_X1   g0951(.A1(new_n1131), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1118), .B2(new_n959), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1130), .A2(new_n1153), .ZN(G378));
  OAI21_X1  g0954(.A(new_n433), .B1(new_n448), .B2(new_n453), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT55), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT55), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1157), .B(new_n433), .C1(new_n448), .C2(new_n453), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n423), .A2(new_n851), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT56), .Z(new_n1160));
  AND3_X1   g0960(.A1(new_n1156), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n916), .B2(G330), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n896), .A2(new_n899), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n911), .A2(new_n910), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n913), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n914), .A2(new_n915), .ZN(new_n1168));
  AND4_X1   g0968(.A1(G330), .A2(new_n1167), .A3(new_n1168), .A4(new_n1163), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n903), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(G330), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1163), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1105), .A2(new_n879), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n902), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n877), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n916), .A2(G330), .A3(new_n1163), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1170), .A2(KEYINPUT122), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1176), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT122), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n1121), .C2(new_n1082), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n690), .A2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1028), .B1(new_n773), .B2(new_n481), .C1(new_n557), .C2(new_n758), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G41), .B(new_n1186), .C1(G68), .C2(new_n777), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n781), .A2(new_n217), .B1(new_n763), .B2(new_n800), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n294), .B(new_n1188), .C1(G283), .C2(new_n795), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(new_n534), .C2(new_n770), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT58), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n202), .B1(new_n255), .B2(G41), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n773), .A2(new_n1146), .B1(new_n776), .B2(new_n415), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n771), .A2(G137), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n1144), .B2(new_n781), .C1(new_n779), .C2(new_n1141), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G125), .C2(new_n786), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT59), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G41), .B1(new_n795), .B2(G124), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G33), .B1(new_n836), .B2(G159), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1191), .A2(new_n1192), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n740), .B1(new_n1201), .B2(new_n749), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(G50), .B2(new_n845), .C1(new_n1172), .C2(new_n751), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT120), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1185), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n959), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1120), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1082), .B1(new_n1118), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1207), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT121), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1178), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n1180), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1178), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1206), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(G375));
  NAND3_X1  g1020(.A1(new_n1091), .A2(new_n1099), .A3(new_n1082), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1127), .A2(new_n986), .A3(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n257), .B1(new_n766), .B2(new_n547), .C1(new_n362), .C2(new_n763), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G294), .A2(new_n786), .B1(new_n788), .B2(G97), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n557), .B2(new_n781), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G283), .C2(new_n774), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1032), .C1(new_n481), .C2(new_n770), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n758), .A2(new_n1144), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n781), .A2(new_n1141), .B1(new_n770), .B2(new_n415), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G137), .C2(new_n774), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n779), .A2(new_n266), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n294), .B1(new_n763), .B2(new_n800), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(G50), .C2(new_n777), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1233), .C1(new_n1146), .C2(new_n766), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n755), .B1(new_n1235), .B2(new_n749), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n873), .B2(new_n751), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n360), .B2(new_n844), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1101), .B2(new_n959), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1222), .A2(new_n1239), .ZN(G381));
  AND2_X1   g1040(.A1(new_n1130), .A2(new_n1153), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1219), .A2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(G381), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G387), .A2(G390), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(G407));
  INV_X1    g1047(.A(G213), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(G343), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1219), .A2(new_n1241), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT123), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(G407), .A2(G213), .A3(new_n1252), .A4(new_n1253), .ZN(G409));
  XNOR2_X1  g1054(.A(G393), .B(G396), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(G390), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n986), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n984), .B2(new_n736), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1006), .B(new_n1007), .C1(new_n1258), .C2(new_n959), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(new_n958), .A3(new_n1078), .A4(new_n1059), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT125), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1255), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1259), .A2(new_n958), .B1(new_n1059), .B2(new_n1078), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1264), .B1(new_n1244), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1255), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1179), .A2(new_n959), .A3(new_n1182), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1205), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n986), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1249), .B1(new_n1274), .B2(new_n1241), .ZN(new_n1275));
  OAI21_X1  g1075(.A(G378), .B1(new_n1206), .B2(new_n1218), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1221), .A2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1091), .A2(new_n1099), .A3(new_n1082), .A4(KEYINPUT60), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(new_n1120), .A3(new_n690), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1239), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n848), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n848), .A2(new_n1282), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1281), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1280), .B2(new_n1239), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1275), .A2(new_n1276), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1275), .A2(new_n1276), .A3(new_n1292), .A4(new_n1288), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1249), .A2(G2897), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1281), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1287), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(G2897), .A3(new_n1249), .A4(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1270), .B1(new_n1294), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1249), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1107), .A2(new_n1110), .A3(new_n1098), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1088), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1208), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1102), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1216), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT121), .B1(new_n1170), .B2(new_n1178), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1310), .B(new_n986), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1205), .A3(new_n1271), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1305), .B1(new_n1314), .B2(G378), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1204), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1317));
  AOI22_X1  g1117(.A1(new_n1316), .A2(new_n1317), .B1(new_n1130), .B2(new_n1153), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1288), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1315), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1321), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1320), .B1(KEYINPUT63), .B2(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT63), .A4(new_n1288), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1269), .B2(new_n1291), .ZN(new_n1326));
  AOI211_X1 g1126(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1263), .C2(new_n1268), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1324), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1323), .A2(new_n1328), .A3(KEYINPUT127), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT127), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1260), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1267), .B1(new_n1266), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1262), .A2(new_n1255), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1291), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT126), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1269), .A2(new_n1325), .A3(new_n1291), .ZN(new_n1336));
  AOI22_X1  g1136(.A1(new_n1320), .A2(KEYINPUT63), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1289), .B1(new_n1303), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1330), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1304), .B1(new_n1329), .B2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(new_n1242), .A2(new_n1276), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1270), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1242), .A2(new_n1276), .A3(new_n1269), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1319), .ZN(G402));
endmodule


