

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743;

  NOR2_X1 U369 ( .A1(G953), .A2(G237), .ZN(n502) );
  XNOR2_X1 U370 ( .A(KEYINPUT3), .B(G119), .ZN(n474) );
  INV_X1 U371 ( .A(G146), .ZN(n460) );
  XNOR2_X1 U372 ( .A(n729), .B(n460), .ZN(n482) );
  BUF_X1 U373 ( .A(n701), .Z(n710) );
  NOR2_X1 U374 ( .A1(n619), .A2(n714), .ZN(n621) );
  NAND2_X2 U375 ( .A1(n388), .A2(n648), .ZN(n584) );
  BUF_X2 U376 ( .A(n664), .Z(n347) );
  XNOR2_X1 U377 ( .A(n535), .B(n534), .ZN(n579) );
  XNOR2_X2 U378 ( .A(n390), .B(n417), .ZN(n459) );
  NOR2_X1 U379 ( .A1(n429), .A2(n560), .ZN(n428) );
  NOR2_X1 U380 ( .A1(n579), .A2(n537), .ZN(n625) );
  INV_X1 U381 ( .A(G953), .ZN(n731) );
  INV_X4 U382 ( .A(G143), .ZN(n458) );
  XNOR2_X1 U383 ( .A(n431), .B(n430), .ZN(n715) );
  NAND2_X1 U384 ( .A1(n428), .A2(n423), .ZN(n431) );
  AND2_X1 U385 ( .A1(n426), .A2(n424), .ZN(n423) );
  NAND2_X1 U386 ( .A1(n387), .A2(n386), .ZN(n385) );
  NOR2_X1 U387 ( .A1(n557), .A2(n518), .ZN(n402) );
  XNOR2_X1 U388 ( .A(n367), .B(KEYINPUT80), .ZN(n634) );
  OR2_X1 U389 ( .A1(n411), .A2(n581), .ZN(n605) );
  XNOR2_X1 U390 ( .A(n691), .B(n690), .ZN(n693) );
  XNOR2_X1 U391 ( .A(n529), .B(n353), .ZN(n575) );
  XOR2_X1 U392 ( .A(n700), .B(KEYINPUT59), .Z(n703) );
  XNOR2_X1 U393 ( .A(n381), .B(n380), .ZN(n551) );
  INV_X1 U394 ( .A(KEYINPUT104), .ZN(n380) );
  NAND2_X1 U395 ( .A1(n384), .A2(n382), .ZN(n381) );
  XNOR2_X1 U396 ( .A(n385), .B(n406), .ZN(n384) );
  NOR2_X2 U397 ( .A1(n372), .A2(G902), .ZN(n535) );
  NOR2_X1 U398 ( .A1(G902), .A2(n712), .ZN(n529) );
  INV_X1 U399 ( .A(KEYINPUT1), .ZN(n421) );
  XNOR2_X1 U400 ( .A(n525), .B(n524), .ZN(n727) );
  OR2_X1 U401 ( .A1(n542), .A2(n407), .ZN(n517) );
  NAND2_X1 U402 ( .A1(n602), .A2(n408), .ZN(n407) );
  INV_X1 U403 ( .A(n531), .ZN(n408) );
  XNOR2_X1 U404 ( .A(n362), .B(KEYINPUT20), .ZN(n526) );
  AND2_X1 U405 ( .A1(n634), .A2(n386), .ZN(n457) );
  INV_X1 U406 ( .A(n576), .ZN(n444) );
  XNOR2_X1 U407 ( .A(G101), .B(G137), .ZN(n478) );
  INV_X1 U408 ( .A(KEYINPUT94), .ZN(n477) );
  XOR2_X1 U409 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n476) );
  INV_X1 U410 ( .A(G134), .ZN(n417) );
  XNOR2_X1 U411 ( .A(G137), .B(KEYINPUT68), .ZN(n524) );
  NOR2_X1 U412 ( .A1(n349), .A2(n425), .ZN(n424) );
  NOR2_X1 U413 ( .A1(n550), .A2(KEYINPUT87), .ZN(n425) );
  AND2_X1 U414 ( .A1(n550), .A2(KEYINPUT87), .ZN(n427) );
  INV_X1 U415 ( .A(KEYINPUT48), .ZN(n413) );
  INV_X1 U416 ( .A(n534), .ZN(n420) );
  XOR2_X1 U417 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n512) );
  XNOR2_X1 U418 ( .A(n404), .B(n508), .ZN(n510) );
  XOR2_X1 U419 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n508) );
  XNOR2_X1 U420 ( .A(n507), .B(n405), .ZN(n404) );
  INV_X1 U421 ( .A(KEYINPUT101), .ZN(n405) );
  XNOR2_X1 U422 ( .A(n365), .B(n501), .ZN(n525) );
  INV_X1 U423 ( .A(G140), .ZN(n441) );
  XNOR2_X1 U424 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n442) );
  INV_X1 U425 ( .A(n585), .ZN(n455) );
  INV_X1 U426 ( .A(n373), .ZN(n599) );
  XNOR2_X1 U427 ( .A(n573), .B(n415), .ZN(n600) );
  XNOR2_X1 U428 ( .A(n574), .B(KEYINPUT39), .ZN(n415) );
  INV_X1 U429 ( .A(KEYINPUT85), .ZN(n574) );
  XNOR2_X1 U430 ( .A(n610), .B(n453), .ZN(n379) );
  INV_X1 U431 ( .A(KEYINPUT111), .ZN(n453) );
  XOR2_X1 U432 ( .A(G478), .B(n516), .Z(n545) );
  INV_X1 U433 ( .A(KEYINPUT28), .ZN(n412) );
  NOR2_X1 U434 ( .A1(n665), .A2(n662), .ZN(n409) );
  XNOR2_X1 U435 ( .A(n359), .B(n473), .ZN(n571) );
  OR2_X1 U436 ( .A1(n530), .A2(n545), .ZN(n373) );
  NAND2_X1 U437 ( .A1(n383), .A2(n398), .ZN(n382) );
  NOR2_X1 U438 ( .A1(n665), .A2(n399), .ZN(n398) );
  XNOR2_X1 U439 ( .A(n402), .B(KEYINPUT86), .ZN(n383) );
  INV_X1 U440 ( .A(KEYINPUT103), .ZN(n406) );
  NAND2_X1 U441 ( .A1(G953), .A2(G902), .ZN(n563) );
  XNOR2_X1 U442 ( .A(n527), .B(KEYINPUT92), .ZN(n528) );
  XNOR2_X1 U443 ( .A(n669), .B(n419), .ZN(n586) );
  INV_X1 U444 ( .A(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U445 ( .A(G116), .B(KEYINPUT9), .ZN(n507) );
  XNOR2_X1 U446 ( .A(n422), .B(KEYINPUT17), .ZN(n488) );
  INV_X1 U447 ( .A(KEYINPUT78), .ZN(n422) );
  XNOR2_X1 U448 ( .A(n460), .B(G125), .ZN(n501) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n495) );
  OR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n493) );
  XNOR2_X1 U451 ( .A(n506), .B(n351), .ZN(n452) );
  XNOR2_X1 U452 ( .A(n578), .B(n577), .ZN(n585) );
  AND2_X1 U453 ( .A1(n575), .A2(n443), .ZN(n578) );
  AND2_X1 U454 ( .A1(n661), .A2(n444), .ZN(n443) );
  NOR2_X1 U455 ( .A1(n545), .A2(n451), .ZN(n602) );
  BUF_X1 U456 ( .A(n586), .Z(n401) );
  XNOR2_X1 U457 ( .A(n482), .B(n483), .ZN(n372) );
  XNOR2_X1 U458 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U459 ( .A(G143), .B(KEYINPUT12), .ZN(n446) );
  XNOR2_X1 U460 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n447) );
  XOR2_X1 U461 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n504) );
  XNOR2_X1 U462 ( .A(n449), .B(n448), .ZN(n375) );
  XNOR2_X1 U463 ( .A(G113), .B(G131), .ZN(n448) );
  XNOR2_X1 U464 ( .A(n450), .B(G104), .ZN(n449) );
  INV_X1 U465 ( .A(G122), .ZN(n450) );
  INV_X1 U466 ( .A(KEYINPUT45), .ZN(n430) );
  AND2_X1 U467 ( .A1(n646), .A2(n369), .ZN(n368) );
  XNOR2_X1 U468 ( .A(n371), .B(n413), .ZN(n370) );
  INV_X1 U469 ( .A(n644), .ZN(n369) );
  AND2_X1 U470 ( .A1(n395), .A2(n572), .ZN(n591) );
  NOR2_X1 U471 ( .A1(n570), .A2(n576), .ZN(n395) );
  NAND2_X1 U472 ( .A1(n545), .A2(n451), .ZN(n592) );
  XNOR2_X1 U473 ( .A(n452), .B(KEYINPUT100), .ZN(n530) );
  XNOR2_X1 U474 ( .A(n727), .B(n363), .ZN(n712) );
  XNOR2_X1 U475 ( .A(n364), .B(n523), .ZN(n363) );
  XNOR2_X1 U476 ( .A(n513), .B(n416), .ZN(n514) );
  XNOR2_X1 U477 ( .A(G107), .B(G122), .ZN(n509) );
  XNOR2_X1 U478 ( .A(n376), .B(n374), .ZN(n700) );
  XNOR2_X1 U479 ( .A(n445), .B(n375), .ZN(n374) );
  XNOR2_X1 U480 ( .A(n525), .B(n505), .ZN(n376) );
  XNOR2_X1 U481 ( .A(n447), .B(n446), .ZN(n445) );
  XNOR2_X1 U482 ( .A(n482), .B(n391), .ZN(n696) );
  XNOR2_X1 U483 ( .A(n471), .B(n463), .ZN(n391) );
  NOR2_X1 U484 ( .A1(G952), .A2(n731), .ZN(n714) );
  XNOR2_X1 U485 ( .A(n437), .B(KEYINPUT42), .ZN(n742) );
  NAND2_X1 U486 ( .A1(n439), .A2(n438), .ZN(n437) );
  INV_X1 U487 ( .A(n605), .ZN(n439) );
  XNOR2_X1 U488 ( .A(n440), .B(n601), .ZN(n743) );
  NAND2_X1 U489 ( .A1(n600), .A2(n599), .ZN(n440) );
  AND2_X1 U490 ( .A1(n377), .A2(n665), .ZN(n642) );
  XNOR2_X1 U491 ( .A(n378), .B(KEYINPUT36), .ZN(n377) );
  NOR2_X1 U492 ( .A1(n379), .A2(n587), .ZN(n378) );
  XNOR2_X1 U493 ( .A(n556), .B(n403), .ZN(n740) );
  XNOR2_X1 U494 ( .A(n555), .B(KEYINPUT32), .ZN(n403) );
  INV_X1 U495 ( .A(KEYINPUT64), .ZN(n555) );
  XNOR2_X1 U496 ( .A(n533), .B(n532), .ZN(n639) );
  NOR2_X1 U497 ( .A1(n605), .A2(n582), .ZN(n367) );
  NOR2_X1 U498 ( .A1(n557), .A2(n393), .ZN(n558) );
  NAND2_X1 U499 ( .A1(n409), .A2(n394), .ZN(n393) );
  INV_X1 U500 ( .A(n579), .ZN(n394) );
  XNOR2_X1 U501 ( .A(n373), .B(KEYINPUT107), .ZN(n636) );
  INV_X1 U502 ( .A(n382), .ZN(n622) );
  XNOR2_X1 U503 ( .A(n571), .B(n421), .ZN(n588) );
  OR2_X1 U504 ( .A1(KEYINPUT47), .A2(n583), .ZN(n348) );
  AND2_X1 U505 ( .A1(n561), .A2(KEYINPUT44), .ZN(n349) );
  INV_X1 U506 ( .A(n662), .ZN(n399) );
  XOR2_X1 U507 ( .A(G131), .B(KEYINPUT4), .Z(n350) );
  XOR2_X1 U508 ( .A(KEYINPUT13), .B(G475), .Z(n351) );
  XOR2_X1 U509 ( .A(KEYINPUT65), .B(n494), .Z(n352) );
  XOR2_X1 U510 ( .A(n528), .B(n456), .Z(n353) );
  XOR2_X1 U511 ( .A(G128), .B(KEYINPUT24), .Z(n354) );
  XOR2_X1 U512 ( .A(KEYINPUT77), .B(KEYINPUT90), .Z(n355) );
  XNOR2_X1 U513 ( .A(n491), .B(KEYINPUT81), .ZN(n356) );
  XOR2_X2 U514 ( .A(G113), .B(G116), .Z(n357) );
  NOR2_X1 U515 ( .A1(n531), .A2(n575), .ZN(n664) );
  XNOR2_X1 U516 ( .A(G122), .B(KEYINPUT16), .ZN(n358) );
  NOR2_X1 U517 ( .A1(n696), .A2(G902), .ZN(n359) );
  NOR2_X1 U518 ( .A1(n599), .A2(n638), .ZN(n654) );
  INV_X1 U519 ( .A(n654), .ZN(n386) );
  AND2_X1 U520 ( .A1(n608), .A2(n609), .ZN(n360) );
  AND2_X1 U521 ( .A1(G224), .A2(n731), .ZN(n361) );
  NAND2_X1 U522 ( .A1(n615), .A2(G234), .ZN(n362) );
  XNOR2_X2 U523 ( .A(KEYINPUT15), .B(G902), .ZN(n615) );
  XNOR2_X1 U524 ( .A(n366), .B(n521), .ZN(n364) );
  XNOR2_X1 U525 ( .A(n520), .B(n354), .ZN(n366) );
  XNOR2_X1 U526 ( .A(n442), .B(n441), .ZN(n365) );
  NAND2_X1 U527 ( .A1(n370), .A2(n368), .ZN(n730) );
  NAND2_X1 U528 ( .A1(n348), .A2(n360), .ZN(n371) );
  XNOR2_X1 U529 ( .A(n372), .B(KEYINPUT112), .ZN(n616) );
  INV_X1 U530 ( .A(n538), .ZN(n387) );
  INV_X1 U531 ( .A(n388), .ZN(n613) );
  XNOR2_X2 U532 ( .A(n492), .B(n356), .ZN(n388) );
  XNOR2_X1 U533 ( .A(n613), .B(KEYINPUT38), .ZN(n649) );
  NAND2_X1 U534 ( .A1(n594), .A2(n388), .ZN(n633) );
  NOR2_X4 U535 ( .A1(n389), .A2(n615), .ZN(n701) );
  NAND2_X1 U536 ( .A1(n686), .A2(n389), .ZN(n687) );
  XNOR2_X2 U537 ( .A(n414), .B(KEYINPUT2), .ZN(n389) );
  XNOR2_X1 U538 ( .A(n390), .B(n355), .ZN(n397) );
  XNOR2_X2 U539 ( .A(n458), .B(G128), .ZN(n390) );
  XNOR2_X1 U540 ( .A(n397), .B(n361), .ZN(n434) );
  XNOR2_X1 U541 ( .A(n436), .B(KEYINPUT46), .ZN(n606) );
  NOR2_X1 U542 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U543 ( .A(n486), .B(n358), .ZN(n432) );
  XNOR2_X1 U544 ( .A(n432), .B(n485), .ZN(n722) );
  OR2_X2 U545 ( .A1(n741), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U546 ( .A1(n392), .A2(n347), .ZN(n418) );
  INV_X1 U547 ( .A(n586), .ZN(n392) );
  NOR2_X2 U548 ( .A1(n546), .A2(n592), .ZN(n549) );
  XNOR2_X2 U549 ( .A(n549), .B(n548), .ZN(n741) );
  NAND2_X1 U550 ( .A1(n701), .A2(G210), .ZN(n692) );
  XNOR2_X1 U551 ( .A(n396), .B(KEYINPUT72), .ZN(n560) );
  NOR2_X2 U552 ( .A1(n559), .A2(n561), .ZN(n396) );
  NOR2_X2 U553 ( .A1(n715), .A2(n730), .ZN(n414) );
  XNOR2_X1 U554 ( .A(n400), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U555 ( .A1(n694), .A2(n714), .ZN(n400) );
  NOR2_X2 U556 ( .A1(n704), .A2(n714), .ZN(n705) );
  XNOR2_X1 U557 ( .A(n580), .B(n412), .ZN(n411) );
  XNOR2_X1 U558 ( .A(n722), .B(n433), .ZN(n689) );
  XNOR2_X1 U559 ( .A(n434), .B(n490), .ZN(n433) );
  INV_X1 U560 ( .A(n675), .ZN(n438) );
  NOR2_X2 U561 ( .A1(n542), .A2(n539), .ZN(n536) );
  NOR2_X1 U562 ( .A1(n588), .A2(n418), .ZN(n541) );
  XNOR2_X2 U563 ( .A(n357), .B(n474), .ZN(n486) );
  NAND2_X1 U564 ( .A1(n410), .A2(KEYINPUT47), .ZN(n589) );
  INV_X1 U565 ( .A(n634), .ZN(n410) );
  NOR2_X1 U566 ( .A1(n581), .A2(n539), .ZN(n572) );
  INV_X1 U567 ( .A(n459), .ZN(n416) );
  XNOR2_X2 U568 ( .A(n535), .B(n420), .ZN(n669) );
  NAND2_X1 U569 ( .A1(n741), .A2(KEYINPUT44), .ZN(n550) );
  NAND2_X1 U570 ( .A1(n551), .A2(n427), .ZN(n426) );
  NOR2_X1 U571 ( .A1(n551), .A2(KEYINPUT87), .ZN(n429) );
  XNOR2_X2 U572 ( .A(n435), .B(n500), .ZN(n542) );
  NOR2_X2 U573 ( .A1(n582), .A2(n499), .ZN(n435) );
  XNOR2_X2 U574 ( .A(n584), .B(n352), .ZN(n582) );
  XNOR2_X2 U575 ( .A(n517), .B(KEYINPUT22), .ZN(n557) );
  NAND2_X1 U576 ( .A1(n743), .A2(n742), .ZN(n436) );
  INV_X1 U577 ( .A(n575), .ZN(n662) );
  INV_X1 U578 ( .A(n452), .ZN(n451) );
  NAND2_X1 U579 ( .A1(n454), .A2(n636), .ZN(n610) );
  NOR2_X1 U580 ( .A1(n401), .A2(n455), .ZN(n454) );
  XOR2_X1 U581 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n456) );
  XNOR2_X1 U582 ( .A(n478), .B(n477), .ZN(n479) );
  INV_X1 U583 ( .A(KEYINPUT69), .ZN(n577) );
  XNOR2_X1 U584 ( .A(n472), .B(G469), .ZN(n473) );
  XNOR2_X1 U585 ( .A(n616), .B(KEYINPUT62), .ZN(n617) );
  XNOR2_X1 U586 ( .A(n515), .B(n514), .ZN(n706) );
  XNOR2_X1 U587 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U588 ( .A(n547), .B(KEYINPUT84), .ZN(n548) );
  INV_X1 U589 ( .A(KEYINPUT63), .ZN(n620) );
  XNOR2_X1 U590 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X2 U591 ( .A(n459), .B(n350), .ZN(n729) );
  XNOR2_X1 U592 ( .A(n524), .B(G140), .ZN(n462) );
  NAND2_X1 U593 ( .A1(G227), .A2(n731), .ZN(n461) );
  XNOR2_X1 U594 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U595 ( .A(G110), .B(G104), .ZN(n469) );
  INV_X1 U596 ( .A(G107), .ZN(n464) );
  NAND2_X1 U597 ( .A1(n464), .A2(KEYINPUT89), .ZN(n467) );
  INV_X1 U598 ( .A(KEYINPUT89), .ZN(n465) );
  NAND2_X1 U599 ( .A1(n465), .A2(G107), .ZN(n466) );
  NAND2_X1 U600 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U601 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U602 ( .A(G101), .B(n470), .ZN(n485) );
  INV_X1 U603 ( .A(n485), .ZN(n471) );
  XNOR2_X1 U604 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n472) );
  INV_X1 U605 ( .A(n588), .ZN(n665) );
  NAND2_X1 U606 ( .A1(n502), .A2(G210), .ZN(n475) );
  XNOR2_X1 U607 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U608 ( .A(n486), .B(n481), .ZN(n483) );
  XNOR2_X1 U609 ( .A(G472), .B(KEYINPUT95), .ZN(n534) );
  INV_X1 U610 ( .A(n401), .ZN(n518) );
  NAND2_X1 U611 ( .A1(G221), .A2(n526), .ZN(n484) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(n484), .Z(n661) );
  XNOR2_X1 U613 ( .A(KEYINPUT93), .B(n661), .ZN(n531) );
  INV_X1 U614 ( .A(KEYINPUT0), .ZN(n500) );
  XNOR2_X1 U615 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n487) );
  XNOR2_X1 U616 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U617 ( .A(n501), .B(n489), .ZN(n490) );
  NAND2_X1 U618 ( .A1(n689), .A2(n615), .ZN(n492) );
  NAND2_X1 U619 ( .A1(G210), .A2(n493), .ZN(n491) );
  NAND2_X1 U620 ( .A1(G214), .A2(n493), .ZN(n648) );
  XOR2_X1 U621 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n494) );
  XNOR2_X1 U622 ( .A(KEYINPUT14), .B(n495), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G952), .A2(n731), .ZN(n566) );
  INV_X1 U624 ( .A(n566), .ZN(n497) );
  NOR2_X1 U625 ( .A1(G898), .A2(n563), .ZN(n496) );
  OR2_X1 U626 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U627 ( .A1(n562), .A2(n498), .ZN(n499) );
  NAND2_X1 U628 ( .A1(G214), .A2(n502), .ZN(n503) );
  XNOR2_X1 U629 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U630 ( .A1(G902), .A2(n700), .ZN(n506) );
  XNOR2_X1 U631 ( .A(n510), .B(n509), .ZN(n515) );
  NAND2_X1 U632 ( .A1(G234), .A2(n731), .ZN(n511) );
  XNOR2_X1 U633 ( .A(n512), .B(n511), .ZN(n522) );
  NAND2_X1 U634 ( .A1(G217), .A2(n522), .ZN(n513) );
  NOR2_X1 U635 ( .A1(G902), .A2(n706), .ZN(n516) );
  XNOR2_X1 U636 ( .A(G119), .B(G110), .ZN(n519) );
  XNOR2_X1 U637 ( .A(n519), .B(KEYINPUT23), .ZN(n521) );
  XOR2_X1 U638 ( .A(KEYINPUT91), .B(KEYINPUT76), .Z(n520) );
  NAND2_X1 U639 ( .A1(n522), .A2(G221), .ZN(n523) );
  NAND2_X1 U640 ( .A1(G217), .A2(n526), .ZN(n527) );
  AND2_X1 U641 ( .A1(n530), .A2(n545), .ZN(n638) );
  INV_X1 U642 ( .A(n347), .ZN(n539) );
  NOR2_X1 U643 ( .A1(n588), .A2(n669), .ZN(n660) );
  NAND2_X1 U644 ( .A1(n536), .A2(n660), .ZN(n533) );
  XNOR2_X1 U645 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n532) );
  NAND2_X1 U646 ( .A1(n536), .A2(n571), .ZN(n537) );
  NOR2_X1 U647 ( .A1(n639), .A2(n625), .ZN(n538) );
  XNOR2_X1 U648 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n540) );
  XNOR2_X1 U649 ( .A(n541), .B(n540), .ZN(n659) );
  NOR2_X1 U650 ( .A1(n659), .A2(n542), .ZN(n544) );
  INV_X1 U651 ( .A(KEYINPUT34), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n544), .B(n543), .ZN(n546) );
  INV_X1 U653 ( .A(KEYINPUT35), .ZN(n547) );
  NAND2_X1 U654 ( .A1(n575), .A2(n401), .ZN(n552) );
  NOR2_X1 U655 ( .A1(n588), .A2(n552), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n553), .B(KEYINPUT79), .ZN(n554) );
  NOR2_X1 U657 ( .A1(n557), .A2(n554), .ZN(n556) );
  XNOR2_X1 U658 ( .A(n558), .B(KEYINPUT105), .ZN(n738) );
  NAND2_X1 U659 ( .A1(n740), .A2(n738), .ZN(n561) );
  INV_X1 U660 ( .A(n562), .ZN(n681) );
  NOR2_X1 U661 ( .A1(n681), .A2(n563), .ZN(n564) );
  XOR2_X1 U662 ( .A(KEYINPUT108), .B(n564), .Z(n565) );
  NOR2_X1 U663 ( .A1(G900), .A2(n565), .ZN(n568) );
  NOR2_X1 U664 ( .A1(n681), .A2(n566), .ZN(n567) );
  NOR2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n579), .A2(n648), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n569), .B(KEYINPUT30), .ZN(n570) );
  INV_X1 U668 ( .A(n571), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n591), .A2(n649), .ZN(n573) );
  AND2_X1 U670 ( .A1(n600), .A2(n638), .ZN(n644) );
  AND2_X1 U671 ( .A1(n579), .A2(n585), .ZN(n580) );
  NOR2_X1 U672 ( .A1(KEYINPUT83), .A2(n457), .ZN(n583) );
  BUF_X1 U673 ( .A(n584), .Z(n587) );
  NOR2_X1 U674 ( .A1(KEYINPUT83), .A2(n589), .ZN(n590) );
  NOR2_X1 U675 ( .A1(n642), .A2(n590), .ZN(n609) );
  NAND2_X1 U676 ( .A1(KEYINPUT83), .A2(n634), .ZN(n598) );
  INV_X1 U677 ( .A(n591), .ZN(n593) );
  NOR2_X1 U678 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U679 ( .A1(KEYINPUT47), .A2(n654), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n633), .A2(n595), .ZN(n596) );
  XOR2_X1 U681 ( .A(KEYINPUT82), .B(n596), .Z(n597) );
  NAND2_X1 U682 ( .A1(n598), .A2(n597), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n601) );
  NAND2_X1 U684 ( .A1(n649), .A2(n648), .ZN(n653) );
  INV_X1 U685 ( .A(n602), .ZN(n651) );
  NOR2_X1 U686 ( .A1(n653), .A2(n651), .ZN(n604) );
  XNOR2_X1 U687 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n604), .B(n603), .ZN(n675) );
  NOR2_X1 U689 ( .A1(n665), .A2(n610), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n611), .A2(n648), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT43), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n646) );
  NAND2_X1 U693 ( .A1(n701), .A2(G472), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(G57) );
  XNOR2_X1 U696 ( .A(n622), .B(G101), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n623), .B(KEYINPUT113), .ZN(G3) );
  NAND2_X1 U698 ( .A1(n625), .A2(n636), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(G104), .ZN(G6) );
  XNOR2_X1 U700 ( .A(G107), .B(KEYINPUT114), .ZN(n629) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n627) );
  NAND2_X1 U702 ( .A1(n625), .A2(n638), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(G9) );
  XOR2_X1 U705 ( .A(G128), .B(KEYINPUT29), .Z(n631) );
  NAND2_X1 U706 ( .A1(n638), .A2(n634), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(G30) );
  XOR2_X1 U708 ( .A(G143), .B(KEYINPUT115), .Z(n632) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n634), .A2(n636), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(G146), .ZN(G48) );
  NAND2_X1 U712 ( .A1(n639), .A2(n636), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(G113), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(KEYINPUT116), .ZN(n641) );
  XNOR2_X1 U716 ( .A(G116), .B(n641), .ZN(G18) );
  XNOR2_X1 U717 ( .A(G125), .B(n642), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n644), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U721 ( .A(G140), .B(KEYINPUT118), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(G42) );
  NOR2_X1 U723 ( .A1(n675), .A2(n659), .ZN(n684) );
  NOR2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U726 ( .A(KEYINPUT119), .B(n652), .Z(n656) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT120), .ZN(n658) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n677) );
  NAND2_X1 U731 ( .A1(n660), .A2(n347), .ZN(n672) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT49), .B(n663), .Z(n668) );
  NOR2_X1 U734 ( .A1(n665), .A2(n347), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(KEYINPUT50), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U739 ( .A(KEYINPUT51), .B(n673), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U742 ( .A(n678), .B(KEYINPUT121), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n679), .B(KEYINPUT52), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n680), .A2(G952), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT122), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n687), .A2(G953), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U750 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n689), .B(KEYINPUT88), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U753 ( .A1(n710), .A2(G469), .ZN(n698) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  NOR2_X1 U755 ( .A1(n714), .A2(n699), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n701), .A2(G475), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U759 ( .A(n706), .B(KEYINPUT123), .Z(n708) );
  NAND2_X1 U760 ( .A1(n710), .A2(G478), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U762 ( .A1(n714), .A2(n709), .ZN(G63) );
  NAND2_X1 U763 ( .A1(G217), .A2(n710), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  NOR2_X1 U766 ( .A1(G953), .A2(n715), .ZN(n720) );
  XOR2_X1 U767 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n717) );
  NAND2_X1 U768 ( .A1(G224), .A2(G953), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(n718) );
  INV_X1 U770 ( .A(G898), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n718), .A2(n721), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n721), .A2(G953), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n724), .B(KEYINPUT125), .ZN(n725) );
  XOR2_X1 U776 ( .A(n726), .B(n725), .Z(G69) );
  XOR2_X1 U777 ( .A(n727), .B(KEYINPUT126), .Z(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n730), .B(n733), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n737) );
  XNOR2_X1 U781 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(G72) );
  XNOR2_X1 U785 ( .A(G110), .B(n738), .ZN(G12) );
  XOR2_X1 U786 ( .A(G119), .B(KEYINPUT127), .Z(n739) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(G21) );
  XOR2_X1 U788 ( .A(n741), .B(G122), .Z(G24) );
  XNOR2_X1 U789 ( .A(n742), .B(G137), .ZN(G39) );
  XNOR2_X1 U790 ( .A(n743), .B(G131), .ZN(G33) );
endmodule

