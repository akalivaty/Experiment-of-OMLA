

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NAND2_X1 U552 ( .A1(G1956), .A2(n736), .ZN(n516) );
  INV_X1 U553 ( .A(KEYINPUT27), .ZN(n698) );
  AND2_X1 U554 ( .A1(n700), .A2(n516), .ZN(n713) );
  INV_X1 U555 ( .A(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U556 ( .A(n719), .B(n718), .ZN(n724) );
  AND2_X1 U557 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U558 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X2 U559 ( .A1(n690), .A2(n794), .ZN(n736) );
  OR2_X1 U560 ( .A1(n689), .A2(n688), .ZN(n793) );
  NOR2_X1 U561 ( .A1(n640), .A2(G651), .ZN(n650) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n538), .Z(n654) );
  NOR2_X1 U563 ( .A1(n526), .A2(n525), .ZN(G164) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n517), .Z(n893) );
  NAND2_X1 U565 ( .A1(G138), .A2(n893), .ZN(n519) );
  INV_X1 U566 ( .A(G2104), .ZN(n521) );
  NOR2_X1 U567 ( .A1(G2105), .A2(n521), .ZN(n896) );
  NAND2_X1 U568 ( .A1(G102), .A2(n896), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n526) );
  AND2_X2 U570 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U571 ( .A1(n889), .A2(G114), .ZN(n520) );
  XNOR2_X1 U572 ( .A(n520), .B(KEYINPUT86), .ZN(n523) );
  AND2_X1 U573 ( .A1(n521), .A2(G2105), .ZN(n888) );
  NAND2_X1 U574 ( .A1(G126), .A2(n888), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT87), .B(n524), .Z(n525) );
  XNOR2_X1 U577 ( .A(G2454), .B(G2443), .ZN(n536) );
  XOR2_X1 U578 ( .A(G2430), .B(KEYINPUT106), .Z(n528) );
  XNOR2_X1 U579 ( .A(G2446), .B(KEYINPUT107), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n528), .B(n527), .ZN(n532) );
  XOR2_X1 U581 ( .A(G2451), .B(G2427), .Z(n530) );
  XNOR2_X1 U582 ( .A(G1348), .B(G1341), .ZN(n529) );
  XNOR2_X1 U583 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U584 ( .A(n532), .B(n531), .Z(n534) );
  XNOR2_X1 U585 ( .A(G2435), .B(G2438), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U587 ( .A(n536), .B(n535), .ZN(n537) );
  AND2_X1 U588 ( .A1(n537), .A2(G14), .ZN(G401) );
  INV_X1 U589 ( .A(G651), .ZN(n541) );
  NOR2_X1 U590 ( .A1(G543), .A2(n541), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G64), .A2(n654), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  NAND2_X1 U593 ( .A1(G52), .A2(n650), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U595 ( .A1(n640), .A2(n541), .ZN(n646) );
  NAND2_X1 U596 ( .A1(G77), .A2(n646), .ZN(n543) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n647) );
  NAND2_X1 U598 ( .A1(G90), .A2(n647), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT9), .B(n544), .ZN(n545) );
  XNOR2_X1 U601 ( .A(KEYINPUT67), .B(n545), .ZN(n546) );
  NOR2_X1 U602 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  NAND2_X1 U605 ( .A1(G101), .A2(n896), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n548), .Z(n551) );
  NAND2_X1 U607 ( .A1(G137), .A2(n893), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT65), .B(n549), .Z(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n689) );
  NAND2_X1 U610 ( .A1(G125), .A2(n888), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G113), .A2(n889), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n687) );
  NOR2_X1 U613 ( .A1(n689), .A2(n687), .ZN(G160) );
  NAND2_X1 U614 ( .A1(G63), .A2(n654), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G51), .A2(n650), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n556), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n647), .A2(G89), .ZN(n557) );
  XNOR2_X1 U619 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U620 ( .A1(G76), .A2(n646), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT5), .B(n560), .Z(n561) );
  XNOR2_X1 U623 ( .A(KEYINPUT72), .B(n561), .ZN(n562) );
  NOR2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(n564), .Z(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n832) );
  NAND2_X1 U630 ( .A1(n832), .A2(G567), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U632 ( .A1(n646), .A2(G68), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT70), .B(n567), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n569) );
  NAND2_X1 U635 ( .A1(G81), .A2(n647), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(n572), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(KEYINPUT68), .Z(n574) );
  NAND2_X1 U640 ( .A1(G56), .A2(n654), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n574), .B(n573), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G43), .A2(n650), .ZN(n575) );
  XNOR2_X1 U643 ( .A(KEYINPUT71), .B(n575), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n985) );
  INV_X1 U646 ( .A(G860), .ZN(n598) );
  OR2_X1 U647 ( .A1(n985), .A2(n598), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G79), .A2(n646), .ZN(n581) );
  NAND2_X1 U651 ( .A1(G92), .A2(n647), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G66), .A2(n654), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G54), .A2(n650), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT15), .B(n586), .Z(n973) );
  OR2_X1 U658 ( .A1(n973), .A2(G868), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G65), .A2(n654), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G53), .A2(n650), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G78), .A2(n646), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G91), .A2(n647), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n970) );
  INV_X1 U667 ( .A(n970), .ZN(G299) );
  INV_X1 U668 ( .A(G868), .ZN(n665) );
  NOR2_X1 U669 ( .A1(G286), .A2(n665), .ZN(n596) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT73), .B(n597), .Z(G297) );
  NAND2_X1 U673 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n599), .A2(n973), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U676 ( .A1(n973), .A2(G868), .ZN(n601) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n601), .ZN(n602) );
  NOR2_X1 U678 ( .A1(G559), .A2(n602), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G868), .A2(n985), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U681 ( .A1(n888), .A2(G123), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G111), .A2(n889), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G135), .A2(n893), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G99), .A2(n896), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n923) );
  XNOR2_X1 U689 ( .A(n923), .B(G2096), .ZN(n613) );
  INV_X1 U690 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G67), .A2(n654), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G55), .A2(n650), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n647), .A2(G93), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT76), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G80), .A2(n646), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U699 ( .A(KEYINPUT77), .B(n619), .Z(n620) );
  OR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n666) );
  NAND2_X1 U701 ( .A1(G559), .A2(n973), .ZN(n622) );
  XOR2_X1 U702 ( .A(n985), .B(n622), .Z(n663) );
  XNOR2_X1 U703 ( .A(KEYINPUT75), .B(n663), .ZN(n623) );
  NOR2_X1 U704 ( .A1(G860), .A2(n623), .ZN(n624) );
  XOR2_X1 U705 ( .A(n666), .B(n624), .Z(G145) );
  NAND2_X1 U706 ( .A1(G72), .A2(n646), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G85), .A2(n647), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT66), .B(n627), .Z(n631) );
  NAND2_X1 U710 ( .A1(G60), .A2(n654), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G47), .A2(n650), .ZN(n628) );
  AND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G48), .A2(n650), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(KEYINPUT78), .ZN(n639) );
  NAND2_X1 U716 ( .A1(G86), .A2(n647), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G61), .A2(n654), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n646), .A2(G73), .ZN(n635) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G49), .A2(n650), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G87), .A2(n640), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U726 ( .A1(n654), .A2(n643), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G651), .A2(G74), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G75), .A2(n646), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G88), .A2(n647), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G50), .A2(n650), .ZN(n651) );
  XNOR2_X1 U733 ( .A(KEYINPUT79), .B(n651), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n654), .A2(G62), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G303) );
  INV_X1 U737 ( .A(G303), .ZN(G166) );
  XOR2_X1 U738 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n657) );
  XNOR2_X1 U739 ( .A(G288), .B(n657), .ZN(n658) );
  XNOR2_X1 U740 ( .A(G305), .B(n658), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n970), .B(G166), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U743 ( .A(n666), .B(n661), .ZN(n662) );
  XNOR2_X1 U744 ( .A(G290), .B(n662), .ZN(n842) );
  XOR2_X1 U745 ( .A(n842), .B(n663), .Z(n664) );
  NOR2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U747 ( .A1(G868), .A2(n666), .ZN(n667) );
  NOR2_X1 U748 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT81), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n672), .B(KEYINPUT21), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n673), .B(KEYINPUT82), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U757 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n676) );
  NAND2_X1 U758 ( .A1(G132), .A2(G82), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U760 ( .A1(n677), .A2(G218), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G96), .A2(n678), .ZN(n840) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n840), .ZN(n679) );
  XNOR2_X1 U763 ( .A(n679), .B(KEYINPUT84), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G108), .A2(G120), .ZN(n680) );
  NOR2_X1 U765 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U766 ( .A1(G69), .A2(n681), .ZN(n841) );
  NAND2_X1 U767 ( .A1(G567), .A2(n841), .ZN(n682) );
  NAND2_X1 U768 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT85), .B(n684), .ZN(G319) );
  INV_X1 U770 ( .A(G319), .ZN(n914) );
  NAND2_X1 U771 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U772 ( .A1(n914), .A2(n685), .ZN(n837) );
  NAND2_X1 U773 ( .A1(n837), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G40), .ZN(n686) );
  OR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  INV_X1 U776 ( .A(n793), .ZN(n690) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U778 ( .A(G1996), .ZN(n943) );
  NOR2_X1 U779 ( .A1(n736), .A2(n943), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n691), .B(KEYINPUT26), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n736), .A2(G1341), .ZN(n693) );
  INV_X1 U782 ( .A(n985), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U785 ( .A(n696), .B(KEYINPUT64), .ZN(n703) );
  NOR2_X1 U786 ( .A1(n973), .A2(n703), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n697), .B(KEYINPUT97), .ZN(n711) );
  INV_X1 U788 ( .A(n736), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n704), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U791 ( .A1(n713), .A2(n970), .ZN(n702) );
  XOR2_X1 U792 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n701) );
  XNOR2_X1 U793 ( .A(n702), .B(n701), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n703), .A2(n973), .ZN(n708) );
  NOR2_X1 U795 ( .A1(n704), .A2(G1348), .ZN(n706) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n736), .ZN(n705) );
  NOR2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U799 ( .A1(n712), .A2(n709), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n717) );
  INV_X1 U801 ( .A(n712), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n713), .A2(n970), .ZN(n714) );
  OR2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n716) );
  AND2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n719) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NOR2_X1 U806 ( .A1(n945), .A2(n736), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT95), .ZN(n722) );
  INV_X1 U808 ( .A(G1961), .ZN(n992) );
  NAND2_X1 U809 ( .A1(n992), .A2(n736), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n729) );
  NAND2_X1 U811 ( .A1(n729), .A2(G171), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n734) );
  NAND2_X1 U813 ( .A1(n736), .A2(G8), .ZN(n773) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n773), .ZN(n748) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n736), .ZN(n745) );
  NOR2_X1 U816 ( .A1(n748), .A2(n745), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT98), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U819 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(n732), .Z(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n746) );
  NAND2_X1 U825 ( .A1(n746), .A2(G286), .ZN(n743) );
  INV_X1 U826 ( .A(G8), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n773), .ZN(n735) );
  XNOR2_X1 U828 ( .A(KEYINPUT99), .B(n735), .ZN(n739) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U830 ( .A1(G166), .A2(n737), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  OR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U833 ( .A(n744), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G8), .A2(n745), .ZN(n750) );
  INV_X1 U835 ( .A(n746), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n770) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n760), .A2(n753), .ZN(n980) );
  XNOR2_X1 U842 ( .A(KEYINPUT100), .B(n980), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n770), .A2(n754), .ZN(n757) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U845 ( .A(n974), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n773), .A2(n755), .ZN(n756) );
  NOR2_X1 U847 ( .A1(KEYINPUT33), .A2(n758), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT101), .ZN(n764) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n967) );
  NAND2_X1 U850 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  OR2_X1 U851 ( .A1(n773), .A2(n761), .ZN(n762) );
  AND2_X1 U852 ( .A1(n967), .A2(n762), .ZN(n763) );
  AND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n769) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U855 ( .A(n765), .B(KEYINPUT94), .Z(n766) );
  XNOR2_X1 U856 ( .A(KEYINPUT24), .B(n766), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n767), .A2(n773), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n776) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n770), .A2(n772), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n811) );
  NAND2_X1 U864 ( .A1(G119), .A2(n888), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G131), .A2(n893), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n896), .A2(G95), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT92), .B(n779), .Z(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n889), .A2(G107), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n874) );
  NAND2_X1 U872 ( .A1(G1991), .A2(n874), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G129), .A2(n888), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G141), .A2(n893), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n896), .A2(G105), .ZN(n786) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n786), .Z(n787) );
  NOR2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n889), .A2(G117), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n875) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n875), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n924) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n825) );
  NAND2_X1 U884 ( .A1(n924), .A2(n825), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(KEYINPUT93), .ZN(n818) );
  INV_X1 U886 ( .A(n818), .ZN(n809) );
  XOR2_X1 U887 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n808) );
  XNOR2_X1 U888 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G128), .A2(n888), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G116), .A2(n889), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U892 ( .A(n799), .B(n798), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G140), .A2(n893), .ZN(n801) );
  NAND2_X1 U894 ( .A1(G104), .A2(n896), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U896 ( .A(KEYINPUT88), .B(n802), .ZN(n803) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n803), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT36), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n808), .B(n807), .ZN(n909) );
  XNOR2_X1 U901 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  NOR2_X1 U902 ( .A1(n909), .A2(n823), .ZN(n934) );
  NAND2_X1 U903 ( .A1(n934), .A2(n825), .ZN(n821) );
  AND2_X1 U904 ( .A1(n809), .A2(n821), .ZN(n810) );
  AND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U907 ( .A1(n982), .A2(n825), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n828) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n875), .ZN(n920) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n874), .ZN(n814) );
  XOR2_X1 U911 ( .A(KEYINPUT103), .B(n814), .Z(n925) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT102), .B(n815), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n925), .A2(n816), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n920), .A2(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n909), .A2(n823), .ZN(n932) );
  NAND2_X1 U920 ( .A1(n824), .A2(n932), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n831) );
  XOR2_X1 U923 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n829) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n829), .ZN(n830) );
  XNOR2_X1 U925 ( .A(n831), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT108), .ZN(G217) );
  NAND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U929 ( .A(G661), .ZN(n834) );
  NOR2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G1), .A2(G3), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n839), .B(KEYINPUT110), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  INV_X1 U937 ( .A(G132), .ZN(G219) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G82), .ZN(G220) );
  NOR2_X1 U941 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XOR2_X1 U943 ( .A(KEYINPUT120), .B(n842), .Z(n844) );
  XNOR2_X1 U944 ( .A(G171), .B(n973), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U946 ( .A(G286), .B(n845), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n846), .B(n985), .ZN(n847) );
  NOR2_X1 U948 ( .A1(G37), .A2(n847), .ZN(G397) );
  XOR2_X1 U949 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2090), .Z(n851) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(G227) );
  XOR2_X1 U958 ( .A(G1981), .B(G1961), .Z(n857) );
  XNOR2_X1 U959 ( .A(G1986), .B(G1966), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n858), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U962 ( .A(G1991), .B(G1996), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U964 ( .A(G2474), .B(G1976), .Z(n862) );
  XNOR2_X1 U965 ( .A(G1956), .B(G1971), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n866) );
  NAND2_X1 U969 ( .A1(G124), .A2(n888), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G112), .A2(n889), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G100), .A2(n896), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n869), .B(KEYINPUT113), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G136), .A2(n893), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U978 ( .A(G162), .B(n874), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n887) );
  NAND2_X1 U980 ( .A1(n896), .A2(G106), .ZN(n877) );
  XOR2_X1 U981 ( .A(KEYINPUT115), .B(n877), .Z(n879) );
  NAND2_X1 U982 ( .A1(n893), .A2(G142), .ZN(n878) );
  NAND2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n880), .B(KEYINPUT45), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G118), .A2(n889), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n888), .A2(G130), .ZN(n883) );
  XOR2_X1 U988 ( .A(KEYINPUT114), .B(n883), .Z(n884) );
  NOR2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U990 ( .A(n887), .B(n886), .Z(n901) );
  NAND2_X1 U991 ( .A1(G127), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G115), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n892), .B(KEYINPUT47), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G139), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G103), .A2(n896), .ZN(n897) );
  XNOR2_X1 U998 ( .A(KEYINPUT117), .B(n897), .ZN(n898) );
  NOR2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n928) );
  XNOR2_X1 U1000 ( .A(G164), .B(n928), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1002 ( .A(KEYINPUT116), .B(KEYINPUT118), .Z(n903) );
  XNOR2_X1 U1003 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G160), .B(n923), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n910), .ZN(n911) );
  XOR2_X1 U1010 ( .A(KEYINPUT119), .B(n911), .Z(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(G397), .A2(n913), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(KEYINPUT121), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(G395), .A2(n916), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n921), .Z(n940) );
  XOR2_X1 U1023 ( .A(G2084), .B(G160), .Z(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n938) );
  XOR2_X1 U1027 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(KEYINPUT50), .B(n931), .ZN(n936) );
  INV_X1 U1031 ( .A(n932), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1038 ( .A(G32), .B(n943), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G27), .B(n945), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(KEYINPUT124), .B(n946), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G1991), .B(G25), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G2072), .B(G33), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT123), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(KEYINPUT53), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G2084), .B(KEYINPUT54), .Z(n957) );
  XNOR2_X1 U1052 ( .A(G34), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(G2090), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G35), .B(n960), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1057 ( .A(KEYINPUT125), .B(n963), .Z(n964) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n964), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n965), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(G11), .ZN(n1019) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT57), .ZN(n989) );
  XNOR2_X1 U1065 ( .A(n970), .B(G1956), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT126), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n1017) );
  INV_X1 U1080 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1081 ( .A(G5), .B(n992), .ZN(n1005) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(G4), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(KEYINPUT127), .B(G1956), .Z(n998) );
  XNOR2_X1 U1089 ( .A(G20), .B(n998), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1001), .Z(n1003) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1095 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

