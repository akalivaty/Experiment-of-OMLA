//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n187), .A2(G107), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n188), .A2(new_n191), .A3(new_n194), .A4(new_n195), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n196), .A2(new_n198), .B1(G101), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n208), .A2(KEYINPUT75), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n206), .B(G146), .C1(new_n202), .C2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n202), .A2(new_n204), .A3(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(KEYINPUT75), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n201), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT10), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT64), .B1(new_n219), .B2(G134), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G137), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n222), .B2(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n219), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n225), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n225), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n188), .A2(new_n191), .A3(new_n195), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT4), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n205), .A2(new_n207), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT0), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n202), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n238), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n212), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n203), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n211), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n201), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n218), .A2(new_n233), .A3(new_n249), .A4(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G140), .ZN(new_n257));
  INV_X1    g071(.A(G953), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(G227), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n257), .B(new_n259), .Z(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n216), .B1(new_n254), .B2(new_n201), .ZN(new_n262));
  INV_X1    g076(.A(new_n233), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n262), .B(new_n263), .C1(KEYINPUT76), .C2(KEYINPUT12), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT12), .B1(new_n263), .B2(KEYINPUT76), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n261), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n218), .A2(new_n249), .A3(new_n255), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n263), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n260), .B1(new_n270), .B2(new_n256), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G469), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n261), .B1(new_n263), .B2(new_n269), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n256), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n264), .B2(new_n267), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(G469), .C1(new_n260), .C2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n275), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G221), .B1(new_n285), .B2(G902), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G214), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n200), .A2(G101), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n236), .B2(new_n237), .ZN(new_n292));
  INV_X1    g106(.A(G119), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G116), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT66), .B(G119), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT5), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G119), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n304), .A3(G113), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(new_n295), .C1(new_n297), .C2(new_n296), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n290), .B1(new_n292), .B2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n201), .A2(KEYINPUT77), .A3(new_n308), .A4(new_n305), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n302), .B2(new_n294), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n238), .A2(new_n313), .A3(new_n248), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G122), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n310), .A2(new_n311), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G224), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT7), .B1(new_n317), .B2(G953), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n244), .B2(new_n246), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n211), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT65), .B1(new_n210), .B2(new_n211), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n324), .A2(new_n325), .A3(new_n208), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n326), .B2(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n322), .B1(new_n254), .B2(new_n321), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n330), .A2(KEYINPUT80), .A3(new_n318), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n292), .A2(new_n309), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n196), .A2(new_n198), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n334), .A2(new_n308), .A3(new_n291), .A4(new_n305), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n315), .B(KEYINPUT8), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT79), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n340), .B(new_n337), .C1(new_n333), .C2(new_n335), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n316), .B(new_n332), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n274), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n315), .A2(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n316), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n317), .A2(G953), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n330), .B(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n345), .A2(new_n355), .A3(new_n358), .A4(new_n356), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n289), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n287), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G472), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n222), .A2(G137), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n219), .A2(G134), .ZN(new_n366));
  OAI21_X1  g180(.A(G131), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n229), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n326), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n205), .A2(new_n207), .B1(new_n241), .B2(new_n242), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n205), .A2(new_n207), .A3(new_n242), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n220), .A2(new_n223), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n227), .A2(new_n228), .ZN(new_n374));
  OAI21_X1  g188(.A(G131), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n372), .B1(new_n375), .B2(new_n229), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n369), .A2(new_n376), .A3(KEYINPUT30), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n247), .B1(new_n230), .B2(new_n232), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n254), .A2(new_n229), .A3(new_n367), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n313), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n308), .A2(new_n312), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G210), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(G101), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT67), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n369), .A2(new_n376), .A3(new_n313), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT30), .B1(new_n369), .B2(new_n376), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n379), .A2(new_n380), .A3(new_n378), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n393), .B1(new_n396), .B2(new_n313), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n383), .A4(new_n390), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n390), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT28), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n313), .B1(new_n369), .B2(new_n376), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n385), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n385), .A2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n406), .A2(new_n383), .B1(new_n397), .B2(new_n390), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n364), .B(new_n274), .C1(new_n400), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n384), .B1(new_n379), .B2(new_n380), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT28), .B1(new_n393), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n385), .A2(new_n402), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT31), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(new_n385), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n401), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n392), .B(new_n399), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n364), .A4(new_n274), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT68), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n411), .A2(new_n390), .A3(new_n412), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n397), .B2(new_n390), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n411), .A2(new_n390), .A3(new_n412), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n420), .B(G472), .C1(new_n428), .C2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n422), .B1(new_n415), .B2(new_n401), .ZN(new_n430));
  INV_X1    g244(.A(new_n427), .ZN(new_n431));
  OAI211_X1 g245(.A(G472), .B(new_n424), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(G472), .A2(G902), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT69), .A3(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n409), .A2(new_n419), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(G125), .A2(G140), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G125), .A2(G140), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT16), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G146), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G140), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n321), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n436), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n204), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT23), .B1(new_n296), .B2(new_n202), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n202), .A2(G119), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n296), .B2(new_n202), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(KEYINPUT23), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G110), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT24), .B(G110), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n441), .B(new_n445), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n448), .A2(new_n452), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT70), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n449), .A2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n439), .A2(new_n440), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n204), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n439), .A2(KEYINPUT71), .A3(G146), .A4(new_n440), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n456), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n454), .A2(new_n464), .A3(new_n468), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n274), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT72), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT25), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT25), .B1(new_n472), .B2(new_n473), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G217), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(G234), .B2(new_n274), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n470), .A2(new_n471), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n478), .A2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT73), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n435), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G122), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G116), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n297), .A2(G122), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G107), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n190), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n202), .A2(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n206), .A2(G128), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n222), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n206), .A3(G128), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  OAI211_X1 g312(.A(G134), .B(new_n497), .C1(new_n498), .C2(new_n496), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n492), .A2(new_n499), .A3(new_n502), .A4(new_n495), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n488), .A2(KEYINPUT14), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n488), .A2(KEYINPUT85), .A3(KEYINPUT14), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n487), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n488), .A2(KEYINPUT14), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n498), .A2(G134), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n495), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n513), .A3(new_n491), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n285), .A2(new_n477), .A3(G953), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n504), .A2(new_n514), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n274), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G478), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n520), .B2(new_n274), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n524), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G475), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n443), .A2(G146), .A3(new_n436), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n445), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n386), .A2(G214), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n206), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n386), .A2(G143), .A3(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n386), .A2(G143), .A3(G214), .ZN(new_n538));
  AOI21_X1  g352(.A(G143), .B1(new_n386), .B2(G214), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n532), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT17), .B(G131), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n225), .A3(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n545), .B2(KEYINPUT17), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n542), .B1(new_n546), .B2(new_n463), .ZN(new_n547));
  XNOR2_X1  g361(.A(G113), .B(G122), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n187), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n549), .B(new_n542), .C1(new_n546), .C2(new_n463), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n530), .B1(new_n553), .B2(new_n274), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n540), .A2(new_n544), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT19), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n444), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n443), .A2(KEYINPUT19), .A3(new_n436), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n204), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n441), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n542), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT82), .A3(new_n550), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n552), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT82), .B1(new_n561), .B2(new_n550), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n530), .B(new_n274), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n550), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n552), .A3(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT20), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n563), .B2(new_n564), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n565), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n554), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G952), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  NAND2_X1  g395(.A1(G234), .A2(G237), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT21), .B(G898), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(G902), .A3(G953), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n529), .A2(new_n579), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n363), .A2(new_n485), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  INV_X1    g406(.A(new_n484), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n274), .B1(new_n400), .B2(new_n407), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n408), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n287), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n589), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n519), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n516), .B1(new_n504), .B2(new_n514), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT33), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n518), .B2(new_n519), .ZN(new_n605));
  OAI211_X1 g419(.A(G478), .B(new_n274), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT33), .B1(new_n601), .B2(new_n602), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n518), .A2(new_n604), .A3(new_n519), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n611), .A2(KEYINPUT89), .A3(G478), .A4(new_n274), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT90), .B(G478), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n521), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n578), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT87), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n361), .A2(new_n618), .A3(new_n288), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n360), .B2(new_n288), .ZN(new_n621));
  AOI211_X1 g435(.A(KEYINPUT88), .B(new_n289), .C1(new_n357), .C2(new_n359), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT81), .B1(new_n342), .B2(new_n274), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n358), .B1(new_n626), .B2(new_n355), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT88), .B1(new_n627), .B2(new_n289), .ZN(new_n628));
  INV_X1    g442(.A(new_n619), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n360), .A2(new_n620), .A3(new_n288), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n617), .B1(new_n623), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n600), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(KEYINPUT92), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT91), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n575), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n565), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n636), .B1(new_n565), .B2(new_n638), .ZN(new_n641));
  OAI22_X1  g455(.A1(new_n640), .A2(new_n641), .B1(new_n637), .B2(new_n575), .ZN(new_n642));
  INV_X1    g456(.A(new_n641), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n637), .A2(new_n575), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n554), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n599), .A3(new_n529), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT93), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n646), .A2(KEYINPUT93), .A3(new_n599), .A4(new_n529), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n623), .A2(new_n631), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n598), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n465), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n482), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n479), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n597), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT94), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n363), .A2(new_n590), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n450), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND2_X1  g480(.A1(new_n623), .A2(new_n631), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n409), .A2(new_n419), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n429), .A2(new_n434), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n287), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n642), .A2(new_n645), .ZN(new_n672));
  INV_X1    g486(.A(new_n554), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n529), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n584), .B1(new_n588), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n667), .A2(new_n671), .A3(new_n658), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n409), .A2(new_n419), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n415), .A2(new_n390), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n403), .A2(new_n385), .A3(new_n401), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n274), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n364), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n681), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n409), .B2(new_n419), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT98), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n360), .A2(new_n361), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT97), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n578), .B1(new_n528), .B2(new_n525), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n288), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n697), .B1(new_n699), .B2(new_n658), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n476), .A2(new_n478), .B1(new_n482), .B2(new_n656), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n698), .A3(KEYINPUT99), .A4(new_n288), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n694), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n692), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n688), .A3(new_n690), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n677), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n287), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n704), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(new_n677), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n616), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n667), .A2(new_n671), .A3(new_n658), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(new_n272), .A2(new_n274), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n286), .A3(new_n275), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n435), .A2(new_n723), .A3(new_n484), .A4(new_n589), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n632), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT101), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n725), .B(new_n727), .ZN(G15));
  NOR3_X1   g542(.A1(new_n435), .A2(new_n723), .A3(new_n484), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n651), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AOI21_X1  g545(.A(new_n701), .B1(new_n623), .B2(new_n631), .ZN(new_n732));
  INV_X1    g546(.A(new_n723), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n670), .A3(new_n590), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND2_X1  g549(.A1(new_n594), .A2(KEYINPUT102), .ZN(new_n736));
  INV_X1    g550(.A(new_n408), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n364), .B1(new_n417), .B2(new_n274), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n594), .A2(KEYINPUT102), .A3(new_n364), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n484), .A3(new_n589), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n667), .A2(new_n742), .A3(new_n698), .A4(new_n733), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n717), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n616), .A2(KEYINPUT103), .A3(new_n716), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n667), .A2(new_n748), .A3(new_n658), .A4(new_n733), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND3_X1  g564(.A1(new_n670), .A2(new_n593), .A3(KEYINPUT104), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n435), .B2(new_n484), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n360), .A2(new_n288), .A3(new_n361), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT103), .B1(new_n616), .B2(new_n716), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n608), .A2(new_n612), .B1(new_n521), .B2(new_n614), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n757), .A2(new_n745), .A3(new_n578), .A4(new_n677), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n287), .B(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT42), .B1(new_n746), .B2(new_n747), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n287), .A2(new_n755), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n485), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n225), .ZN(G33));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n485), .A3(new_n678), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n279), .A2(new_n260), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n276), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n277), .B(KEYINPUT45), .C1(new_n260), .C2(new_n279), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(G469), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n771), .A3(new_n774), .A4(G469), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n281), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n275), .B1(new_n776), .B2(KEYINPUT46), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n286), .B(new_n710), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n613), .A2(new_n615), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n578), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT43), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n785), .A3(new_n578), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n658), .A2(new_n596), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT106), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT106), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n658), .A2(new_n790), .A3(new_n596), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT44), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(KEYINPUT44), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n781), .A2(new_n755), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  INV_X1    g610(.A(new_n755), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n286), .B1(new_n778), .B2(new_n779), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT47), .B(new_n286), .C1(new_n778), .C2(new_n779), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n670), .A2(new_n593), .A3(new_n717), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NOR3_X1   g619(.A1(new_n797), .A2(new_n583), .A3(new_n723), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n691), .A3(new_n593), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n617), .ZN(new_n808));
  INV_X1    g622(.A(new_n754), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n784), .A2(new_n584), .A3(new_n786), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n723), .A3(new_n797), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n810), .A2(new_n484), .A3(new_n741), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n667), .A3(new_n733), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n581), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n658), .A3(new_n739), .A4(new_n740), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n782), .A2(new_n579), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n807), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n814), .A2(new_n289), .A3(new_n695), .A4(new_n733), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT50), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(KEYINPUT50), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n822), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n800), .A2(new_n801), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g645(.A(new_n722), .ZN(new_n832));
  INV_X1    g646(.A(new_n275), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(new_n286), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n800), .A2(new_n837), .A3(new_n801), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n814), .A2(new_n755), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n829), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n821), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n826), .B2(new_n828), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n800), .A2(new_n801), .A3(new_n836), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(new_n840), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT51), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g662(.A(new_n808), .B(new_n816), .C1(new_n843), .C2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n734), .A2(new_n725), .A3(new_n730), .A4(new_n743), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT107), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n651), .A2(new_n729), .B1(new_n632), .B2(new_n724), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(KEYINPUT107), .A3(new_n734), .A4(new_n743), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n663), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n617), .B1(new_n675), .B2(new_n579), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n600), .A2(new_n362), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n859), .A3(new_n591), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n435), .A2(new_n674), .A3(new_n529), .A4(new_n677), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n658), .B(new_n762), .C1(new_n748), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n766), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n863), .B2(new_n766), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n865), .A2(new_n866), .A3(new_n764), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n861), .A3(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n689), .A2(new_n658), .A3(new_n677), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n667), .A2(new_n287), .A3(new_n698), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n679), .A2(new_n719), .A3(new_n749), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT52), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n850), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n766), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT108), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n760), .A2(new_n763), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n863), .A2(new_n864), .A3(new_n766), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n860), .A3(new_n851), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n871), .A2(KEYINPUT109), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n871), .A2(KEYINPUT109), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT111), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n873), .A2(new_n886), .A3(KEYINPUT111), .A4(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n860), .B1(new_n853), .B2(new_n855), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n883), .A2(new_n893), .A3(new_n867), .A4(new_n885), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n894), .A2(KEYINPUT110), .A3(new_n850), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT110), .B1(new_n894), .B2(new_n850), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n868), .A2(new_n850), .A3(new_n872), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n849), .B(new_n892), .C1(new_n898), .C2(new_n887), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n580), .A2(new_n258), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n593), .B(new_n286), .C1(new_n835), .C2(KEYINPUT49), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n706), .B(new_n902), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n903));
  INV_X1    g717(.A(new_n783), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n288), .A3(new_n691), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(G75));
  XOR2_X1   g720(.A(new_n352), .B(KEYINPUT115), .Z(new_n907));
  XOR2_X1   g721(.A(new_n354), .B(KEYINPUT55), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(G210), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n913), .B(new_n274), .C1(new_n873), .C2(new_n886), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n914), .B2(KEYINPUT56), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n258), .A2(G952), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n873), .A2(new_n886), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G210), .A3(G902), .ZN(new_n919));
  INV_X1    g733(.A(new_n912), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n911), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT117), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n915), .A2(new_n924), .A3(new_n921), .A4(new_n917), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n918), .B(new_n887), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n281), .B(KEYINPUT57), .Z(new_n928));
  OAI21_X1  g742(.A(new_n272), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n274), .B1(new_n873), .B2(new_n886), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(new_n775), .A3(new_n773), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n916), .B1(new_n929), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  INV_X1    g747(.A(new_n570), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n916), .ZN(G60));
  XNOR2_X1  g751(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n611), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n917), .B1(new_n927), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n892), .B1(new_n898), .B2(new_n887), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  INV_X1    g759(.A(new_n611), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n873), .B2(new_n886), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n656), .B(KEYINPUT119), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n917), .C1(new_n480), .C2(new_n950), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  NOR2_X1   g769(.A1(new_n893), .A2(G953), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n258), .B1(new_n585), .B2(G224), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(new_n907), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(G898), .B2(new_n258), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  NAND4_X1  g777(.A1(new_n781), .A2(new_n667), .A3(new_n698), .A4(new_n809), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n876), .A2(new_n766), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n802), .B2(new_n803), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n275), .A3(new_n777), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n793), .A3(new_n286), .A4(new_n710), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n755), .B1(new_n792), .B2(KEYINPUT44), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n749), .A2(new_n679), .A3(new_n719), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT124), .B1(new_n795), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n964), .B(new_n966), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n795), .A2(KEYINPUT124), .A3(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n981), .A2(new_n982), .A3(new_n964), .A4(new_n966), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n978), .A2(new_n258), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n396), .B(KEYINPUT121), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n557), .A2(new_n558), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n258), .B1(G227), .B2(G900), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n987), .B(KEYINPUT122), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n711), .A2(new_n797), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n485), .A3(new_n858), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n969), .B2(new_n970), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n795), .A2(KEYINPUT123), .A3(new_n994), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n975), .A2(new_n714), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n975), .A2(new_n714), .A3(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n999), .A2(new_n1004), .A3(new_n804), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n992), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n989), .A2(new_n991), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G72));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n999), .A2(new_n1004), .A3(new_n804), .A4(new_n893), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n433), .B(KEYINPUT63), .Z(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n683), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g829(.A(KEYINPUT127), .B(new_n683), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n917), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n397), .A2(new_n401), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n978), .A2(new_n893), .A3(new_n983), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n1012), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n898), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1022), .A2(new_n683), .A3(new_n1012), .A4(new_n1018), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1021), .A2(new_n1023), .ZN(G57));
endmodule


