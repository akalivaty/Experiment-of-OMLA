

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745;

  XNOR2_X1 U377 ( .A(n397), .B(n396), .ZN(n458) );
  AND2_X1 U378 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U379 ( .A1(G902), .A2(n705), .ZN(n475) );
  XNOR2_X1 U380 ( .A(n395), .B(G119), .ZN(n407) );
  OR2_X1 U381 ( .A1(n537), .A2(n523), .ZN(n554) );
  XNOR2_X1 U382 ( .A(n541), .B(n540), .ZN(n617) );
  OR2_X2 U383 ( .A1(n530), .A2(n651), .ZN(n533) );
  XNOR2_X2 U384 ( .A(n527), .B(KEYINPUT32), .ZN(n543) );
  XNOR2_X2 U385 ( .A(n514), .B(KEYINPUT102), .ZN(n542) );
  INV_X2 U386 ( .A(G953), .ZN(n649) );
  NOR2_X1 U387 ( .A1(n732), .A2(KEYINPUT81), .ZN(n401) );
  AND2_X1 U388 ( .A1(n617), .A2(n544), .ZN(n375) );
  XNOR2_X1 U389 ( .A(n579), .B(KEYINPUT106), .ZN(n745) );
  XNOR2_X1 U390 ( .A(n554), .B(n386), .ZN(n637) );
  AND2_X1 U391 ( .A1(n561), .A2(n528), .ZN(n549) );
  XNOR2_X1 U392 ( .A(n477), .B(G125), .ZN(n437) );
  INV_X2 U393 ( .A(KEYINPUT68), .ZN(n415) );
  INV_X2 U394 ( .A(KEYINPUT69), .ZN(n365) );
  XNOR2_X1 U395 ( .A(n599), .B(KEYINPUT82), .ZN(n732) );
  OR2_X2 U396 ( .A1(n693), .A2(n597), .ZN(n424) );
  XNOR2_X2 U397 ( .A(n484), .B(n409), .ZN(n719) );
  XNOR2_X1 U398 ( .A(n437), .B(n436), .ZN(n724) );
  INV_X1 U399 ( .A(KEYINPUT10), .ZN(n436) );
  XNOR2_X1 U400 ( .A(n729), .B(n417), .ZN(n478) );
  INV_X1 U401 ( .A(KEYINPUT0), .ZN(n396) );
  XNOR2_X1 U402 ( .A(G113), .B(KEYINPUT71), .ZN(n406) );
  XNOR2_X1 U403 ( .A(n466), .B(G137), .ZN(n491) );
  NAND2_X1 U404 ( .A1(n379), .A2(n400), .ZN(n378) );
  INV_X1 U405 ( .A(KEYINPUT2), .ZN(n400) );
  XNOR2_X1 U406 ( .A(n424), .B(n423), .ZN(n511) );
  XNOR2_X1 U407 ( .A(n384), .B(n383), .ZN(n465) );
  INV_X1 U408 ( .A(KEYINPUT8), .ZN(n383) );
  XNOR2_X1 U409 ( .A(n724), .B(n462), .ZN(n463) );
  XNOR2_X1 U410 ( .A(G128), .B(G119), .ZN(n460) );
  XOR2_X1 U411 ( .A(KEYINPUT93), .B(G110), .Z(n461) );
  XNOR2_X1 U412 ( .A(G116), .B(G107), .ZN(n445) );
  XOR2_X1 U413 ( .A(KEYINPUT7), .B(G122), .Z(n446) );
  XNOR2_X1 U414 ( .A(n441), .B(n440), .ZN(n604) );
  XNOR2_X1 U415 ( .A(n724), .B(n403), .ZN(n440) );
  XNOR2_X1 U416 ( .A(n478), .B(n420), .ZN(n496) );
  OR2_X1 U417 ( .A1(n668), .A2(n562), .ZN(n563) );
  XNOR2_X1 U418 ( .A(n426), .B(n376), .ZN(n580) );
  INV_X1 U419 ( .A(KEYINPUT19), .ZN(n376) );
  AND2_X1 U420 ( .A1(n511), .A2(n669), .ZN(n426) );
  XNOR2_X1 U421 ( .A(n366), .B(KEYINPUT28), .ZN(n583) );
  NOR2_X1 U422 ( .A1(n560), .A2(n561), .ZN(n366) );
  INV_X1 U423 ( .A(KEYINPUT95), .ZN(n394) );
  INV_X1 U424 ( .A(KEYINPUT22), .ZN(n399) );
  XNOR2_X1 U425 ( .A(KEYINPUT16), .B(G122), .ZN(n408) );
  XOR2_X1 U426 ( .A(G122), .B(G104), .Z(n432) );
  XOR2_X1 U427 ( .A(G143), .B(G113), .Z(n434) );
  XNOR2_X1 U428 ( .A(n476), .B(G134), .ZN(n727) );
  INV_X1 U429 ( .A(KEYINPUT45), .ZN(n372) );
  NAND2_X1 U430 ( .A1(n367), .A2(n595), .ZN(n599) );
  XNOR2_X1 U431 ( .A(n368), .B(n592), .ZN(n367) );
  XNOR2_X1 U432 ( .A(G107), .B(G104), .ZN(n419) );
  XNOR2_X1 U433 ( .A(KEYINPUT77), .B(G110), .ZN(n418) );
  XNOR2_X1 U434 ( .A(n727), .B(G146), .ZN(n494) );
  XNOR2_X1 U435 ( .A(n491), .B(n490), .ZN(n725) );
  NAND2_X1 U436 ( .A1(G237), .A2(G234), .ZN(n430) );
  AND2_X1 U437 ( .A1(n508), .A2(n637), .ZN(n571) );
  AND2_X1 U438 ( .A1(n529), .A2(n404), .ZN(n508) );
  XNOR2_X1 U439 ( .A(n443), .B(n442), .ZN(n537) );
  XNOR2_X1 U440 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U441 ( .A(n382), .B(n444), .ZN(n451) );
  BUF_X1 U442 ( .A(n692), .Z(n704) );
  XNOR2_X1 U443 ( .A(n412), .B(n411), .ZN(n413) );
  AND2_X1 U444 ( .A1(n607), .A2(G953), .ZN(n710) );
  XNOR2_X1 U445 ( .A(n389), .B(n387), .ZN(n644) );
  XNOR2_X1 U446 ( .A(n388), .B(KEYINPUT98), .ZN(n387) );
  NAND2_X1 U447 ( .A1(n371), .A2(n660), .ZN(n389) );
  INV_X1 U448 ( .A(KEYINPUT31), .ZN(n388) );
  AND2_X1 U449 ( .A1(n582), .A2(n583), .ZN(n638) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n626) );
  INV_X1 U451 ( .A(KEYINPUT97), .ZN(n390) );
  OR2_X1 U452 ( .A1(n632), .A2(n589), .ZN(n356) );
  INV_X1 U453 ( .A(G146), .ZN(n477) );
  NOR2_X1 U454 ( .A1(n598), .A2(n732), .ZN(n357) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(G137), .Z(n358) );
  XOR2_X1 U456 ( .A(n586), .B(KEYINPUT80), .Z(n359) );
  AND2_X1 U457 ( .A1(n553), .A2(n552), .ZN(n360) );
  AND2_X1 U458 ( .A1(n501), .A2(n651), .ZN(n361) );
  AND2_X1 U459 ( .A1(n572), .A2(n526), .ZN(n362) );
  NOR2_X1 U460 ( .A1(n513), .A2(n654), .ZN(n363) );
  AND2_X1 U461 ( .A1(n431), .A2(n507), .ZN(n364) );
  BUF_X1 U462 ( .A(n515), .Z(n654) );
  XNOR2_X2 U463 ( .A(n365), .B(G131), .ZN(n476) );
  NAND2_X1 U464 ( .A1(n638), .A2(n665), .ZN(n584) );
  NAND2_X1 U465 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U466 ( .A(n568), .B(n567), .ZN(n369) );
  NOR2_X1 U467 ( .A1(n591), .A2(n590), .ZN(n370) );
  XNOR2_X1 U468 ( .A(n496), .B(n495), .ZN(n620) );
  AND2_X1 U469 ( .A1(n405), .A2(n561), .ZN(n520) );
  XNOR2_X2 U470 ( .A(n563), .B(KEYINPUT41), .ZN(n685) );
  INV_X1 U471 ( .A(n547), .ZN(n371) );
  NAND2_X1 U472 ( .A1(n580), .A2(n364), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n486), .B(n485), .ZN(n611) );
  NAND2_X1 U474 ( .A1(n378), .A2(n597), .ZN(n377) );
  NAND2_X1 U475 ( .A1(n371), .A2(n686), .ZN(n535) );
  XNOR2_X2 U476 ( .A(n373), .B(n372), .ZN(n598) );
  NAND2_X1 U477 ( .A1(n360), .A2(n374), .ZN(n373) );
  XNOR2_X1 U478 ( .A(n375), .B(KEYINPUT44), .ZN(n374) );
  AND2_X2 U479 ( .A1(n380), .A2(n377), .ZN(n603) );
  NAND2_X1 U480 ( .A1(n401), .A2(n402), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n381), .A2(KEYINPUT81), .ZN(n380) );
  NAND2_X1 U482 ( .A1(n357), .A2(n597), .ZN(n381) );
  NAND2_X1 U483 ( .A1(n465), .A2(G217), .ZN(n382) );
  NAND2_X1 U484 ( .A1(n649), .A2(G234), .ZN(n384) );
  XNOR2_X1 U485 ( .A(n385), .B(KEYINPUT36), .ZN(n573) );
  AND2_X1 U486 ( .A1(n570), .A2(n571), .ZN(n385) );
  INV_X1 U487 ( .A(KEYINPUT104), .ZN(n386) );
  NAND2_X1 U488 ( .A1(n626), .A2(n644), .ZN(n551) );
  NAND2_X1 U489 ( .A1(n393), .A2(n392), .ZN(n391) );
  INV_X1 U490 ( .A(n654), .ZN(n392) );
  XNOR2_X1 U491 ( .A(n548), .B(n394), .ZN(n393) );
  XNOR2_X2 U492 ( .A(G116), .B(KEYINPUT3), .ZN(n395) );
  INV_X1 U493 ( .A(n458), .ZN(n547) );
  NAND2_X1 U494 ( .A1(n398), .A2(n363), .ZN(n514) );
  NAND2_X1 U495 ( .A1(n398), .A2(n362), .ZN(n527) );
  NAND2_X1 U496 ( .A1(n398), .A2(n361), .ZN(n552) );
  XNOR2_X2 U497 ( .A(n459), .B(n399), .ZN(n398) );
  INV_X1 U498 ( .A(n598), .ZN(n402) );
  XNOR2_X2 U499 ( .A(n475), .B(n474), .ZN(n561) );
  XNOR2_X2 U500 ( .A(n575), .B(KEYINPUT38), .ZN(n668) );
  BUF_X2 U501 ( .A(n511), .Z(n575) );
  XNOR2_X2 U502 ( .A(n447), .B(n416), .ZN(n729) );
  XNOR2_X2 U503 ( .A(n415), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U505 ( .A(n439), .B(n438), .Z(n403) );
  AND2_X1 U506 ( .A1(n559), .A2(n669), .ZN(n404) );
  NOR2_X1 U507 ( .A1(n518), .A2(n545), .ZN(n405) );
  XNOR2_X1 U508 ( .A(n410), .B(KEYINPUT88), .ZN(n412) );
  XNOR2_X1 U509 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n462) );
  XNOR2_X1 U510 ( .A(n494), .B(n478), .ZN(n486) );
  XNOR2_X1 U511 ( .A(n705), .B(n706), .ZN(n707) );
  XNOR2_X1 U512 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X2 U513 ( .A(n407), .B(n406), .ZN(n484) );
  XNOR2_X1 U514 ( .A(n408), .B(KEYINPUT74), .ZN(n409) );
  XNOR2_X1 U515 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n410) );
  NAND2_X1 U516 ( .A1(n649), .A2(G224), .ZN(n411) );
  XNOR2_X1 U517 ( .A(n413), .B(n437), .ZN(n414) );
  XNOR2_X1 U518 ( .A(n719), .B(n414), .ZN(n421) );
  XNOR2_X2 U519 ( .A(G143), .B(G128), .ZN(n447) );
  XNOR2_X1 U520 ( .A(KEYINPUT66), .B(G101), .ZN(n417) );
  XNOR2_X1 U521 ( .A(n419), .B(n418), .ZN(n717) );
  XNOR2_X1 U522 ( .A(n717), .B(KEYINPUT72), .ZN(n420) );
  XNOR2_X1 U523 ( .A(n421), .B(n496), .ZN(n693) );
  XNOR2_X1 U524 ( .A(KEYINPUT15), .B(G902), .ZN(n596) );
  INV_X1 U525 ( .A(n596), .ZN(n597) );
  INV_X1 U526 ( .A(G902), .ZN(n487) );
  INV_X1 U527 ( .A(G237), .ZN(n422) );
  NAND2_X1 U528 ( .A1(n487), .A2(n422), .ZN(n425) );
  AND2_X1 U529 ( .A1(n425), .A2(G210), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n425), .A2(G214), .ZN(n669) );
  XNOR2_X1 U531 ( .A(G898), .B(KEYINPUT89), .ZN(n714) );
  NAND2_X1 U532 ( .A1(n714), .A2(G953), .ZN(n427) );
  XOR2_X1 U533 ( .A(KEYINPUT90), .B(n427), .Z(n720) );
  NAND2_X1 U534 ( .A1(n720), .A2(G902), .ZN(n428) );
  NAND2_X1 U535 ( .A1(n649), .A2(G952), .ZN(n504) );
  NAND2_X1 U536 ( .A1(n428), .A2(n504), .ZN(n431) );
  INV_X1 U537 ( .A(KEYINPUT14), .ZN(n429) );
  XNOR2_X1 U538 ( .A(n430), .B(n429), .ZN(n683) );
  INV_X1 U539 ( .A(n683), .ZN(n507) );
  XNOR2_X1 U540 ( .A(n476), .B(G140), .ZN(n433) );
  XNOR2_X1 U541 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U542 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U543 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n439) );
  NOR2_X1 U544 ( .A1(G953), .A2(G237), .ZN(n480) );
  NAND2_X1 U545 ( .A1(G214), .A2(n480), .ZN(n438) );
  NAND2_X1 U546 ( .A1(n604), .A2(n487), .ZN(n443) );
  XNOR2_X1 U547 ( .A(KEYINPUT13), .B(G475), .ZN(n442) );
  XNOR2_X1 U548 ( .A(KEYINPUT100), .B(G478), .ZN(n453) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n444) );
  XNOR2_X1 U550 ( .A(n446), .B(n445), .ZN(n449) );
  XOR2_X1 U551 ( .A(G134), .B(n447), .Z(n448) );
  XNOR2_X1 U552 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n701) );
  NOR2_X1 U554 ( .A1(G902), .A2(n701), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n453), .B(n452), .ZN(n536) );
  AND2_X1 U556 ( .A1(n537), .A2(n536), .ZN(n671) );
  NAND2_X1 U557 ( .A1(n596), .A2(G234), .ZN(n454) );
  XNOR2_X1 U558 ( .A(n454), .B(KEYINPUT20), .ZN(n471) );
  AND2_X1 U559 ( .A1(n471), .A2(G221), .ZN(n456) );
  INV_X1 U560 ( .A(KEYINPUT21), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n456), .B(n455), .ZN(n655) );
  INV_X1 U562 ( .A(n655), .ZN(n528) );
  AND2_X1 U563 ( .A1(n671), .A2(n528), .ZN(n457) );
  NAND2_X1 U564 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U565 ( .A(n461), .B(n460), .ZN(n464) );
  XOR2_X1 U566 ( .A(n464), .B(n463), .Z(n470) );
  NAND2_X1 U567 ( .A1(G221), .A2(n465), .ZN(n468) );
  INV_X1 U568 ( .A(G140), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n491), .B(KEYINPUT24), .ZN(n467) );
  XNOR2_X1 U570 ( .A(n470), .B(n469), .ZN(n705) );
  XOR2_X1 U571 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n473) );
  NAND2_X1 U572 ( .A1(n471), .A2(G217), .ZN(n472) );
  XOR2_X1 U573 ( .A(n473), .B(n472), .Z(n474) );
  INV_X1 U574 ( .A(n561), .ZN(n519) );
  XNOR2_X1 U575 ( .A(KEYINPUT96), .B(KEYINPUT76), .ZN(n479) );
  XNOR2_X1 U576 ( .A(n358), .B(n479), .ZN(n482) );
  NAND2_X1 U577 ( .A1(n480), .A2(G210), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U579 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U580 ( .A1(n611), .A2(n487), .ZN(n488) );
  XNOR2_X2 U581 ( .A(n488), .B(G472), .ZN(n515) );
  INV_X1 U582 ( .A(KEYINPUT6), .ZN(n489) );
  XNOR2_X2 U583 ( .A(n515), .B(n489), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n519), .A2(n529), .ZN(n501) );
  INV_X1 U585 ( .A(KEYINPUT91), .ZN(n490) );
  NAND2_X1 U586 ( .A1(n649), .A2(G227), .ZN(n492) );
  XNOR2_X1 U587 ( .A(n725), .B(n492), .ZN(n493) );
  OR2_X2 U588 ( .A1(n620), .A2(G902), .ZN(n498) );
  XNOR2_X1 U589 ( .A(KEYINPUT70), .B(G469), .ZN(n497) );
  XNOR2_X2 U590 ( .A(n498), .B(n497), .ZN(n581) );
  INV_X1 U591 ( .A(KEYINPUT64), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n499), .B(KEYINPUT1), .ZN(n500) );
  XNOR2_X1 U593 ( .A(n581), .B(n500), .ZN(n651) );
  XNOR2_X1 U594 ( .A(G101), .B(KEYINPUT110), .ZN(n502) );
  XNOR2_X1 U595 ( .A(n552), .B(n502), .ZN(G3) );
  NAND2_X1 U596 ( .A1(n519), .A2(n651), .ZN(n513) );
  INV_X1 U597 ( .A(n513), .ZN(n509) );
  INV_X1 U598 ( .A(n536), .ZN(n523) );
  NOR2_X1 U599 ( .A1(G900), .A2(n649), .ZN(n503) );
  NAND2_X1 U600 ( .A1(n503), .A2(G902), .ZN(n505) );
  NAND2_X1 U601 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U602 ( .A1(n507), .A2(n506), .ZN(n518) );
  NOR2_X1 U603 ( .A1(n655), .A2(n518), .ZN(n559) );
  NAND2_X1 U604 ( .A1(n509), .A2(n571), .ZN(n510) );
  XNOR2_X1 U605 ( .A(n510), .B(KEYINPUT43), .ZN(n512) );
  INV_X1 U606 ( .A(n575), .ZN(n569) );
  NAND2_X1 U607 ( .A1(n512), .A2(n569), .ZN(n593) );
  XNOR2_X1 U608 ( .A(n593), .B(G140), .ZN(G42) );
  XNOR2_X1 U609 ( .A(n542), .B(G110), .ZN(G12) );
  AND2_X1 U610 ( .A1(n515), .A2(n669), .ZN(n517) );
  XOR2_X1 U611 ( .A(KEYINPUT105), .B(KEYINPUT30), .Z(n516) );
  XNOR2_X1 U612 ( .A(n517), .B(n516), .ZN(n521) );
  NAND2_X1 U613 ( .A1(n528), .A2(n581), .ZN(n545) );
  NAND2_X1 U614 ( .A1(n521), .A2(n520), .ZN(n578) );
  NOR2_X1 U615 ( .A1(n578), .A2(n668), .ZN(n522) );
  XNOR2_X1 U616 ( .A(n522), .B(KEYINPUT39), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n537), .A2(n523), .ZN(n525) );
  INV_X1 U618 ( .A(KEYINPUT101), .ZN(n524) );
  XNOR2_X1 U619 ( .A(n525), .B(n524), .ZN(n643) );
  OR2_X1 U620 ( .A1(n555), .A2(n643), .ZN(n594) );
  XNOR2_X1 U621 ( .A(n594), .B(G134), .ZN(G36) );
  XNOR2_X1 U622 ( .A(n651), .B(KEYINPUT87), .ZN(n572) );
  NOR2_X1 U623 ( .A1(n529), .A2(n561), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n543), .B(G119), .ZN(G21) );
  NAND2_X1 U625 ( .A1(n549), .A2(n529), .ZN(n530) );
  INV_X1 U626 ( .A(KEYINPUT73), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n531), .B(KEYINPUT33), .ZN(n532) );
  XNOR2_X2 U628 ( .A(n533), .B(n532), .ZN(n686) );
  INV_X1 U629 ( .A(KEYINPUT34), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n535), .B(n534), .ZN(n539) );
  OR2_X1 U631 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n538), .B(KEYINPUT103), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n539), .A2(n576), .ZN(n541) );
  INV_X1 U634 ( .A(KEYINPUT35), .ZN(n540) );
  OR2_X1 U635 ( .A1(n519), .A2(n545), .ZN(n546) );
  NOR2_X1 U636 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U637 ( .A1(n549), .A2(n654), .ZN(n550) );
  NOR2_X1 U638 ( .A1(n550), .A2(n651), .ZN(n660) );
  NAND2_X1 U639 ( .A1(n643), .A2(n554), .ZN(n665) );
  NAND2_X1 U640 ( .A1(n551), .A2(n665), .ZN(n553) );
  OR2_X2 U641 ( .A1(n555), .A2(n554), .ZN(n558) );
  XNOR2_X1 U642 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n556) );
  XNOR2_X1 U643 ( .A(n556), .B(KEYINPUT107), .ZN(n557) );
  XNOR2_X1 U644 ( .A(n558), .B(n557), .ZN(n618) );
  NAND2_X1 U645 ( .A1(n654), .A2(n559), .ZN(n560) );
  AND2_X1 U646 ( .A1(n583), .A2(n581), .ZN(n564) );
  NAND2_X1 U647 ( .A1(n671), .A2(n669), .ZN(n562) );
  NAND2_X1 U648 ( .A1(n564), .A2(n685), .ZN(n566) );
  INV_X1 U649 ( .A(KEYINPUT42), .ZN(n565) );
  XNOR2_X1 U650 ( .A(n566), .B(n565), .ZN(n744) );
  NOR2_X1 U651 ( .A1(n618), .A2(n744), .ZN(n568) );
  XOR2_X1 U652 ( .A(KEYINPUT83), .B(KEYINPUT46), .Z(n567) );
  NOR2_X1 U653 ( .A1(n561), .A2(n569), .ZN(n570) );
  NAND2_X1 U654 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X2 U655 ( .A(n574), .B(KEYINPUT109), .ZN(n742) );
  XNOR2_X1 U656 ( .A(n742), .B(KEYINPUT84), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n579) );
  AND2_X1 U659 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n584), .A2(KEYINPUT47), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n745), .A2(n585), .ZN(n586) );
  INV_X1 U662 ( .A(n638), .ZN(n632) );
  XNOR2_X1 U663 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n587), .A2(n665), .ZN(n588) );
  XOR2_X1 U665 ( .A(KEYINPUT75), .B(n588), .Z(n589) );
  NAND2_X1 U666 ( .A1(n359), .A2(n356), .ZN(n590) );
  INV_X1 U667 ( .A(KEYINPUT48), .ZN(n592) );
  AND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U669 ( .A(n599), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n598), .A2(n601), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT78), .ZN(n647) );
  NOR2_X2 U673 ( .A1(n603), .A2(n647), .ZN(n692) );
  NAND2_X1 U674 ( .A1(n692), .A2(G475), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT59), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n606), .B(n605), .ZN(n608) );
  INV_X1 U677 ( .A(G952), .ZN(n607) );
  NOR2_X2 U678 ( .A1(n608), .A2(n710), .ZN(n610) );
  XOR2_X1 U679 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n609) );
  XNOR2_X1 U680 ( .A(n610), .B(n609), .ZN(G60) );
  NAND2_X1 U681 ( .A1(n692), .A2(G472), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT62), .B(n611), .Z(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U684 ( .A1(n614), .A2(n710), .ZN(n616) );
  XNOR2_X1 U685 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n616), .B(n615), .ZN(G57) );
  XNOR2_X1 U687 ( .A(n617), .B(G122), .ZN(G24) );
  XOR2_X1 U688 ( .A(n618), .B(G131), .Z(G33) );
  NAND2_X1 U689 ( .A1(n704), .A2(G469), .ZN(n622) );
  XOR2_X1 U690 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n619) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n623), .A2(n710), .ZN(G54) );
  INV_X1 U694 ( .A(n637), .ZN(n641) );
  NOR2_X1 U695 ( .A1(n641), .A2(n626), .ZN(n625) );
  XNOR2_X1 U696 ( .A(G104), .B(KEYINPUT111), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(G6) );
  NOR2_X1 U698 ( .A1(n643), .A2(n626), .ZN(n631) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n628) );
  XNOR2_X1 U700 ( .A(G107), .B(KEYINPUT112), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(KEYINPUT26), .B(n629), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n631), .B(n630), .ZN(G9) );
  NOR2_X1 U704 ( .A1(n632), .A2(n643), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n634) );
  XNOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G30) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT116), .ZN(n640) );
  XNOR2_X1 U711 ( .A(G146), .B(n640), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n641), .A2(n644), .ZN(n642) );
  XOR2_X1 U713 ( .A(G113), .B(n642), .Z(G15) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U715 ( .A(G116), .B(n645), .Z(G18) );
  NOR2_X1 U716 ( .A1(n357), .A2(KEYINPUT2), .ZN(n646) );
  XOR2_X1 U717 ( .A(KEYINPUT79), .B(n646), .Z(n648) );
  OR2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n690) );
  INV_X1 U720 ( .A(n651), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n652), .A2(n549), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT50), .ZN(n659) );
  AND2_X1 U723 ( .A1(n519), .A2(n655), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n656), .B(KEYINPUT49), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n392), .A2(n657), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n661) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n662), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n663), .A2(n685), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT117), .B(n664), .ZN(n680) );
  NAND2_X1 U731 ( .A1(n665), .A2(n669), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n666), .A2(n668), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT118), .ZN(n675) );
  INV_X1 U734 ( .A(n668), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n673) );
  INV_X1 U736 ( .A(n671), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U739 ( .A(n686), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT119), .B(n678), .Z(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U745 ( .A1(n684), .A2(G952), .ZN(n688) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n691), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n692), .A2(G210), .ZN(n698) );
  XOR2_X1 U751 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U752 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n693), .B(n696), .ZN(n697) );
  XNOR2_X1 U755 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X2 U756 ( .A1(n699), .A2(n710), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n700), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U758 ( .A1(n704), .A2(G478), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U760 ( .A1(n710), .A2(n703), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n704), .A2(G217), .ZN(n708) );
  XOR2_X1 U762 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n706) );
  NOR2_X1 U763 ( .A1(n710), .A2(n709), .ZN(G66) );
  NOR2_X1 U764 ( .A1(n598), .A2(G953), .ZN(n711) );
  XOR2_X1 U765 ( .A(KEYINPUT123), .B(n711), .Z(n716) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n712) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(n712), .Z(n713) );
  NOR2_X1 U768 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n723) );
  XNOR2_X1 U770 ( .A(n717), .B(G101), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n719), .B(n718), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U773 ( .A(n723), .B(n722), .Z(G69) );
  XOR2_X1 U774 ( .A(n725), .B(n724), .Z(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U776 ( .A(n728), .B(KEYINPUT124), .Z(n731) );
  XNOR2_X1 U777 ( .A(n729), .B(KEYINPUT125), .ZN(n730) );
  XNOR2_X1 U778 ( .A(n731), .B(n730), .ZN(n735) );
  BUF_X1 U779 ( .A(n732), .Z(n733) );
  XOR2_X1 U780 ( .A(n735), .B(n733), .Z(n734) );
  NOR2_X1 U781 ( .A1(n734), .A2(G953), .ZN(n740) );
  XNOR2_X1 U782 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G953), .ZN(n738) );
  XOR2_X1 U785 ( .A(KEYINPUT126), .B(n738), .Z(n739) );
  NOR2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U787 ( .A(KEYINPUT127), .B(n741), .ZN(G72) );
  XNOR2_X1 U788 ( .A(n742), .B(G125), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U790 ( .A(G137), .B(n744), .Z(G39) );
  XNOR2_X1 U791 ( .A(G143), .B(n745), .ZN(G45) );
endmodule

