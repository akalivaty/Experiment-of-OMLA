//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n202), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT65), .B(G244), .Z(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G77), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n212), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n226), .B(new_n229), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT13), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n253), .B(G274), .C1(G41), .C2(G45), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT66), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G226), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G232), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT67), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n257), .B(new_n260), .C1(new_n264), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G97), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n266), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n255), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n223), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n252), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n270), .B2(new_n273), .ZN(new_n284));
  NOR4_X1   g0084(.A1(new_n284), .A2(KEYINPUT13), .A3(new_n281), .A4(new_n255), .ZN(new_n285));
  OAI21_X1  g0085(.A(G169), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n283), .A2(new_n285), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G179), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n254), .B(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n268), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n259), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n272), .B1(new_n294), .B2(new_n257), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n282), .B(new_n291), .C1(new_n295), .C2(new_n276), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT13), .ZN(new_n297));
  AOI211_X1 g0097(.A(new_n256), .B(new_n259), .C1(new_n292), .C2(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n277), .B1(new_n298), .B2(new_n272), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(new_n252), .A3(new_n282), .A4(new_n291), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT14), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n302), .A3(G169), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n287), .A2(new_n289), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G20), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n266), .A2(G20), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(KEYINPUT76), .B1(new_n307), .B2(G77), .ZN(new_n308));
  INV_X1    g0108(.A(G20), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n308), .B1(KEYINPUT76), .B2(new_n306), .C1(new_n309), .C2(G68), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT69), .B1(new_n206), .B2(new_n266), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n312), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n230), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT11), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n253), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n222), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n309), .A2(G1), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n322), .A2(new_n325), .A3(new_n314), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G68), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n316), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n304), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n288), .A2(G190), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n331), .C1(new_n332), .C2(new_n288), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n321), .A2(new_n219), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT73), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n326), .A2(G77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n219), .A2(G20), .ZN(new_n337));
  OR2_X1    g0137(.A1(KEYINPUT8), .A2(G58), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT8), .A2(G58), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n305), .A3(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n337), .A2(KEYINPUT72), .A3(new_n340), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT15), .B(G87), .Z(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n309), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT72), .B1(new_n337), .B2(new_n340), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n341), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n311), .A2(new_n230), .A3(new_n313), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n335), .B(new_n336), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G179), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n218), .A2(new_n276), .A3(new_n279), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n291), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT71), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n291), .A2(KEYINPUT71), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G1698), .B1(new_n264), .B2(new_n269), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n292), .A2(new_n293), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT68), .A3(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(G238), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n361), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G107), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(G232), .A3(new_n258), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n357), .B1(new_n367), .B2(new_n277), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n350), .B1(new_n351), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(G169), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n330), .A2(new_n333), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n338), .A2(new_n339), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n307), .B1(G20), .B2(new_n203), .ZN(new_n375));
  INV_X1    g0175(.A(G150), .ZN(new_n376));
  INV_X1    g0176(.A(new_n305), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n314), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n326), .A2(G50), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n380), .C1(G50), .C2(new_n321), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n360), .A2(G223), .A3(new_n362), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n361), .A2(G222), .A3(new_n258), .ZN(new_n383));
  INV_X1    g0183(.A(new_n219), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n361), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n255), .B1(new_n385), .B2(new_n277), .ZN(new_n386));
  INV_X1    g0186(.A(new_n280), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G226), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n381), .B1(new_n389), .B2(G179), .ZN(new_n390));
  INV_X1    g0190(.A(G169), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n389), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(G190), .A3(new_n388), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n381), .B(KEYINPUT9), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n386), .A2(new_n388), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n332), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n332), .B1(new_n386), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT10), .B1(new_n398), .B2(KEYINPUT75), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n398), .A2(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n401), .A3(KEYINPUT10), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n267), .A2(new_n309), .A3(new_n268), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n309), .A4(new_n268), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n407), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n411), .A3(G68), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n207), .A2(new_n222), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n305), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n292), .A2(new_n293), .A3(new_n309), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n405), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n408), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n416), .B1(new_n421), .B2(G68), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n314), .B(new_n418), .C1(new_n422), .C2(KEYINPUT16), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n321), .A2(new_n373), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n326), .B2(new_n373), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n213), .A2(G1698), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n428), .C1(new_n261), .C2(new_n262), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n276), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n255), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n391), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n431), .A2(new_n255), .A3(new_n433), .A4(new_n351), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT18), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n440), .B(new_n437), .C1(new_n423), .C2(new_n425), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n425), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT77), .B1(new_n404), .B2(new_n405), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n410), .B1(new_n408), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n416), .B1(new_n445), .B2(G68), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n348), .B1(new_n446), .B2(KEYINPUT16), .ZN(new_n447));
  INV_X1    g0247(.A(new_n408), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n419), .B2(new_n405), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n417), .B1(new_n449), .B2(new_n222), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT16), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n443), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n432), .A2(new_n434), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G200), .ZN(new_n455));
  INV_X1    g0255(.A(new_n454), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT78), .A2(G190), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT78), .A2(G190), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n453), .A2(KEYINPUT17), .A3(new_n455), .A4(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n423), .A2(new_n425), .A3(new_n455), .A4(new_n461), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT17), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n442), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n350), .B1(new_n368), .B2(new_n332), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT74), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n368), .A2(G190), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n350), .B(KEYINPUT74), .C1(new_n368), .C2(new_n332), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n372), .A2(new_n403), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n292), .A2(new_n293), .A3(G303), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n267), .A2(new_n268), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n215), .A2(G1698), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n477), .B(new_n478), .C1(G257), .C2(G1698), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n276), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(G274), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n484), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n487), .A2(G270), .A3(new_n276), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n309), .C1(G33), .C2(new_n271), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n314), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n314), .A2(KEYINPUT20), .A3(new_n493), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n322), .A2(new_n492), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n253), .A2(G33), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n348), .A2(G116), .A3(new_n321), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n491), .B(new_n505), .C1(new_n459), .C2(new_n490), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n490), .A3(G169), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(new_n490), .A3(KEYINPUT21), .A4(G169), .ZN(new_n510));
  INV_X1    g0310(.A(new_n486), .ZN(new_n511));
  NOR4_X1   g0311(.A1(new_n480), .A2(new_n351), .A3(new_n511), .A4(new_n488), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n509), .A3(new_n510), .A4(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n322), .A2(new_n271), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n348), .A2(new_n321), .A3(new_n502), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n271), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n305), .A2(G77), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n271), .A2(new_n214), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G20), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n519), .B(new_n525), .C1(new_n449), .C2(new_n214), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n518), .B1(new_n526), .B2(new_n314), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  INV_X1    g0329(.A(G244), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT4), .B1(new_n267), .B2(new_n268), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n258), .B(new_n531), .C1(new_n532), .C2(new_n530), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n292), .A2(new_n293), .B1(new_n210), .B2(G1698), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n529), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n494), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n277), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n487), .A2(new_n276), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n511), .B1(new_n538), .B2(G257), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n351), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n276), .B1(new_n535), .B2(new_n494), .ZN(new_n541));
  INV_X1    g0341(.A(new_n539), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n391), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n528), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n537), .A2(new_n539), .ZN(new_n546));
  INV_X1    g0346(.A(G190), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n527), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n223), .A2(new_n258), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n530), .A2(G1698), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n261), .C2(new_n262), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n276), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n253), .A2(G45), .ZN(new_n556));
  AND2_X1   g0356(.A1(G33), .A2(G41), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(G250), .C1(new_n557), .C2(new_n230), .ZN(new_n558));
  INV_X1    g0358(.A(G274), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n556), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n209), .A2(new_n271), .A3(new_n214), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT19), .B(new_n563), .C1(new_n272), .C2(G20), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n309), .B(G68), .C1(new_n261), .C2(new_n262), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n344), .B2(new_n271), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n314), .B1(new_n322), .B2(new_n343), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n348), .A2(G87), .A3(new_n321), .A4(new_n502), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n555), .B2(new_n560), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n562), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n314), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n348), .A2(new_n321), .A3(new_n342), .A4(new_n502), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n322), .A2(new_n343), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n561), .A2(new_n351), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n391), .B1(new_n555), .B2(new_n560), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n554), .A2(G20), .ZN(new_n582));
  OAI211_X1 g0382(.A(KEYINPUT22), .B(new_n309), .C1(new_n261), .C2(new_n262), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(G87), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  OAI211_X1 g0386(.A(G20), .B(new_n214), .C1(new_n586), .C2(KEYINPUT79), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(KEYINPUT79), .ZN(new_n588));
  XOR2_X1   g0388(.A(new_n587), .B(new_n588), .Z(new_n589));
  AOI211_X1 g0389(.A(G20), .B(new_n209), .C1(new_n292), .C2(new_n293), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n585), .B(new_n589), .C1(new_n590), .C2(KEYINPUT22), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT24), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n361), .A2(new_n309), .A3(G87), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n589), .A4(new_n585), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n348), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n321), .A2(new_n599), .A3(G107), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT25), .B1(new_n322), .B2(new_n214), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n600), .A2(new_n601), .B1(new_n214), .B2(new_n517), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n210), .A2(new_n258), .ZN(new_n604));
  OAI221_X1 g0404(.A(new_n604), .B1(G257), .B2(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n277), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n538), .A2(G264), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n609), .A3(new_n486), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n332), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(G190), .B2(new_n610), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n581), .B1(new_n603), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n391), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n610), .A2(G179), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n598), .C2(new_n602), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n515), .A2(new_n550), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n475), .A2(new_n617), .ZN(G372));
  AND2_X1   g0418(.A1(new_n400), .A2(new_n402), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n426), .B2(new_n438), .ZN(new_n622));
  AOI211_X1 g0422(.A(KEYINPUT82), .B(new_n437), .C1(new_n423), .C2(new_n425), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n440), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT82), .B1(new_n453), .B2(new_n437), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n426), .A2(new_n621), .A3(new_n438), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(KEYINPUT18), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n333), .A2(new_n370), .A3(new_n369), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(new_n330), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n466), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n392), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n616), .A2(new_n509), .A3(new_n510), .A4(new_n513), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n569), .A2(new_n574), .B1(new_n561), .B2(new_n351), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT80), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n555), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n555), .A2(new_n635), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n560), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n638), .B2(G169), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n544), .A2(new_n548), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n573), .A2(new_n575), .A3(new_n570), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT81), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT81), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n569), .A2(new_n643), .A3(new_n570), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n562), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n636), .A2(new_n637), .ZN(new_n646));
  INV_X1    g0446(.A(new_n560), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n332), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n603), .B2(new_n612), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n633), .A2(new_n640), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n647), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G200), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(new_n562), .A3(new_n642), .A4(new_n644), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n527), .B1(new_n546), .B2(new_n391), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n540), .A4(new_n639), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT26), .ZN(new_n657));
  INV_X1    g0457(.A(new_n639), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n580), .A2(new_n528), .A3(new_n540), .A4(new_n543), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n651), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n632), .B1(new_n475), .B2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(new_n616), .ZN(new_n664));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n253), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n603), .A2(new_n673), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n603), .B2(new_n612), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n664), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n509), .A2(new_n510), .A3(new_n513), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n673), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n674), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n504), .A2(new_n672), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT83), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n514), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n677), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n682), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n227), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n563), .A2(G116), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n234), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n661), .A2(new_n673), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT87), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n544), .A2(new_n548), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n700), .A2(new_n633), .A3(new_n650), .A4(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n639), .B1(new_n645), .B2(new_n648), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n544), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n658), .B1(new_n706), .B2(KEYINPUT86), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n659), .A2(new_n705), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT86), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n709), .C1(new_n656), .C2(new_n705), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n699), .B1(new_n711), .B2(new_n673), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n698), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n514), .A2(new_n549), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n613), .A3(new_n616), .A4(new_n673), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n638), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n546), .A3(new_n610), .A4(new_n490), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n541), .A2(new_n542), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n561), .A2(new_n608), .A3(new_n609), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n537), .A2(new_n512), .A3(new_n539), .A4(new_n719), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT84), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT84), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n718), .A2(new_n725), .A3(new_n512), .A4(new_n719), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(KEYINPUT85), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT85), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n723), .A2(new_n732), .A3(new_n726), .A4(new_n724), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n721), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n734), .B2(new_n672), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n713), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT88), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n696), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR3_X1   g0540(.A1(new_n309), .A2(new_n351), .A3(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n460), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G322), .ZN(new_n743));
  INV_X1    g0543(.A(G311), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n547), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n309), .A2(new_n351), .A3(new_n332), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G190), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n459), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n361), .B1(new_n752), .B2(G326), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n332), .A2(G179), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G20), .A3(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G20), .A3(new_n547), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n756), .A2(G303), .B1(new_n759), .B2(G329), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n751), .A2(new_n753), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n754), .A2(G20), .A3(new_n547), .ZN(new_n763));
  INV_X1    g0563(.A(G294), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n309), .B1(new_n757), .B2(G190), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n761), .B1(new_n762), .B2(new_n763), .C1(new_n764), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(G87), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n361), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT91), .Z(new_n772));
  INV_X1    g0572(.A(new_n763), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  INV_X1    g0574(.A(new_n742), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G58), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n752), .B1(new_n749), .B2(G68), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n772), .A2(new_n774), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n768), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G97), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n758), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n780), .B(new_n783), .C1(new_n384), .C2(new_n745), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n769), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n231), .B1(new_n309), .B2(G169), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT90), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n693), .B1(G45), .B2(new_n666), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n361), .A2(G355), .A3(new_n227), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G116), .B2(new_n227), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT89), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n690), .A2(new_n477), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n233), .A2(new_n482), .A3(G50), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n247), .B2(new_n482), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n788), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n791), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n802), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n789), .B(new_n804), .C1(new_n686), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n687), .A2(new_n791), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n686), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n371), .A2(new_n672), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n349), .A2(new_n672), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n473), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n812), .B2(new_n371), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n697), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(new_n737), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n791), .ZN(new_n816));
  INV_X1    g0616(.A(new_n745), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n752), .A2(G303), .B1(new_n817), .B2(G116), .ZN(new_n818));
  INV_X1    g0618(.A(new_n749), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n762), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT93), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n759), .A2(G311), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n763), .A2(new_n209), .B1(new_n755), .B2(new_n214), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n361), .B(new_n823), .C1(G294), .C2(new_n775), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n821), .A2(new_n780), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n775), .A2(G143), .B1(new_n752), .B2(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n376), .B2(new_n819), .C1(new_n781), .C2(new_n745), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n477), .B1(new_n755), .B2(new_n202), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G132), .B2(new_n759), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n828), .B(new_n830), .C1(new_n207), .C2(new_n768), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n763), .A2(new_n222), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n825), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G77), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n788), .A2(new_n800), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n833), .A2(new_n788), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n836), .B(new_n790), .C1(new_n813), .C2(new_n801), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n816), .A2(new_n837), .ZN(G384));
  OAI21_X1  g0638(.A(new_n474), .B1(new_n712), .B2(new_n698), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n632), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n329), .A2(new_n672), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n302), .B1(new_n301), .B2(G169), .ZN(new_n843));
  AOI211_X1 g0643(.A(KEYINPUT14), .B(new_n391), .C1(new_n297), .C2(new_n300), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n283), .A2(new_n285), .A3(new_n351), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n333), .B(new_n842), .C1(new_n846), .C2(new_n328), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n328), .A2(new_n673), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n304), .A2(KEYINPUT94), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT94), .B1(new_n304), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT95), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT95), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n847), .B(new_n853), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n670), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n447), .B1(KEYINPUT16), .B2(new_n446), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n425), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(new_n442), .C2(new_n466), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n857), .A2(new_n425), .B1(new_n437), .B2(new_n670), .ZN(new_n860));
  INV_X1    g0660(.A(new_n463), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n426), .A2(new_n438), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n426), .A2(new_n856), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n463), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n812), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n661), .A2(new_n873), .A3(new_n371), .A4(new_n673), .ZN(new_n874));
  INV_X1    g0674(.A(new_n810), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n855), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT96), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n624), .A2(new_n627), .A3(new_n670), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  INV_X1    g0681(.A(new_n466), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n864), .B1(new_n628), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n866), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n463), .B(new_n864), .C1(new_n622), .C2(new_n623), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n869), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT39), .B1(new_n887), .B2(new_n871), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n870), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n304), .A2(new_n329), .A3(new_n673), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n880), .A2(new_n881), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n841), .B(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n813), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n852), .B2(new_n854), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n896), .A2(new_n715), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n734), .A2(new_n672), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT31), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT97), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT97), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n901), .B(KEYINPUT31), .C1(new_n734), .C2(new_n672), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n897), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n887), .B2(new_n871), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(new_n855), .A3(new_n872), .A4(new_n813), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n904), .A2(new_n906), .B1(new_n907), .B2(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n474), .A2(new_n903), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(G330), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n893), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n253), .B2(new_n666), .ZN(new_n913));
  OAI211_X1 g0713(.A(G20), .B(new_n231), .C1(new_n524), .C2(KEYINPUT35), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n492), .B(new_n914), .C1(KEYINPUT35), .C2(new_n524), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI21_X1  g0716(.A(new_n219), .B1(new_n207), .B2(new_n222), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n917), .A2(new_n234), .B1(G50), .B2(new_n222), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n665), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n752), .A2(G143), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n202), .B2(new_n745), .C1(new_n819), .C2(new_n781), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n361), .B1(new_n742), .B2(new_n376), .ZN(new_n923));
  INV_X1    g0723(.A(G137), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n755), .A2(new_n207), .B1(new_n924), .B2(new_n758), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n926), .B1(new_n222), .B2(new_n768), .C1(new_n384), .C2(new_n763), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n773), .A2(G97), .ZN(new_n928));
  INV_X1    g0728(.A(new_n752), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n928), .B1(new_n819), .B2(new_n764), .C1(new_n929), .C2(new_n744), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n477), .B(new_n930), .C1(G317), .C2(new_n759), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n755), .A2(new_n492), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT46), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT101), .Z(new_n934));
  OAI22_X1  g0734(.A1(new_n932), .A2(KEYINPUT46), .B1(new_n762), .B2(new_n745), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n779), .B2(G107), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(G303), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n742), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n927), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n791), .B1(new_n942), .B2(new_n788), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n803), .B1(new_n227), .B2(new_n343), .C1(new_n243), .C2(new_n796), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n673), .B1(new_n642), .B2(new_n644), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n658), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n704), .B2(new_n945), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n943), .B(new_n944), .C1(new_n805), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n666), .A2(G45), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(G1), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n700), .B(new_n702), .C1(new_n527), .C2(new_n673), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n655), .A2(new_n540), .A3(new_n672), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n951), .A2(KEYINPUT99), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT99), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n682), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT45), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n682), .A2(new_n955), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n688), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT100), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n681), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n687), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n677), .A2(new_n680), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n739), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n739), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n691), .B(KEYINPUT41), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n950), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n955), .A2(new_n681), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT42), .Z(new_n975));
  INV_X1    g0775(.A(new_n955), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n664), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n672), .B1(new_n977), .B2(new_n544), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n973), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n688), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n948), .B1(new_n972), .B2(new_n983), .ZN(G387));
  NAND2_X1  g0784(.A1(new_n374), .A2(new_n202), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n694), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n482), .C1(KEYINPUT50), .C2(new_n985), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G68), .B2(G77), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n795), .B1(new_n240), .B2(new_n482), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n361), .A2(new_n227), .A3(new_n694), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n227), .A2(G107), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n803), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n749), .A2(G311), .B1(new_n817), .B2(G303), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT104), .B(G322), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n994), .B1(new_n995), .B2(new_n742), .C1(new_n929), .C2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(new_n1000), .B1(G283), .B2(new_n779), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n764), .B2(new_n755), .C1(new_n1000), .C2(new_n999), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT49), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n759), .A2(G326), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n477), .B1(new_n773), .B2(G116), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n768), .A2(new_n343), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n929), .A2(new_n781), .B1(new_n222), .B2(new_n745), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n374), .C2(new_n749), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n756), .A2(new_n219), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n759), .A2(G150), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n928), .A2(new_n1012), .A3(new_n477), .A4(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT103), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1011), .B(new_n1015), .C1(new_n202), .C2(new_n742), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n993), .B1(new_n1017), .B2(new_n787), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n791), .B(new_n1018), .C1(new_n677), .C2(new_n802), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n966), .B2(new_n950), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n691), .B(KEYINPUT106), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n967), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n966), .A2(new_n739), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(G393));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n961), .B2(new_n968), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n961), .B2(new_n968), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n955), .A2(new_n802), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n803), .B1(new_n271), .B2(new_n227), .C1(new_n250), .C2(new_n796), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n774), .B1(new_n762), .B2(new_n755), .C1(new_n758), .C2(new_n997), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n364), .B1(new_n764), .B2(new_n745), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n492), .B2(new_n768), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n775), .A2(G311), .B1(new_n752), .B2(G317), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT107), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1035), .B2(KEYINPUT52), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(KEYINPUT52), .B2(new_n1035), .C1(new_n938), .C2(new_n819), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n929), .A2(new_n376), .B1(new_n781), .B2(new_n742), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT51), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n779), .A2(G77), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n749), .A2(G50), .B1(new_n817), .B2(new_n374), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n477), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n773), .B2(G87), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n759), .A2(G143), .ZN(new_n1044));
  AND4_X1   g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1039), .B(new_n1045), .C1(new_n222), .C2(new_n755), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n791), .B1(new_n1047), .B2(new_n788), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1028), .A2(new_n1029), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n961), .B2(new_n950), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1027), .A2(new_n1050), .ZN(G390));
  OAI211_X1 g0851(.A(new_n813), .B(G330), .C1(new_n730), .C2(new_n735), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n854), .A3(new_n852), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT109), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT109), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1055), .A3(new_n854), .A4(new_n852), .ZN(new_n1056));
  INV_X1    g0856(.A(G330), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n894), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n903), .A2(new_n855), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n876), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1052), .B1(new_n854), .B2(new_n852), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n812), .A2(new_n371), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n711), .A2(new_n673), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n875), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n903), .A2(new_n1058), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1063), .B(new_n1067), .C1(new_n1068), .C2(new_n855), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n839), .B(new_n632), .C1(new_n1057), .C2(new_n909), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n854), .A2(new_n852), .B1(new_n874), .B2(new_n875), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n890), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n888), .A2(new_n889), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n855), .A2(new_n1066), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n887), .B2(new_n871), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT108), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1062), .B(new_n1076), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1059), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n888), .A2(new_n889), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n622), .A2(new_n623), .A3(new_n440), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT18), .B1(new_n625), .B2(new_n626), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n882), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n864), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n885), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n866), .B1(new_n1092), .B2(new_n865), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT38), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n871), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n890), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n854), .A2(new_n852), .B1(new_n1065), .B2(new_n875), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT108), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1085), .A2(new_n1086), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1073), .B(new_n1082), .C1(new_n1083), .C2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1071), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1082), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1083), .B1(new_n1104), .B2(new_n1076), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(new_n1022), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n929), .A2(new_n1108), .B1(new_n745), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G132), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n819), .A2(new_n924), .B1(new_n1112), .B2(new_n742), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n756), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT53), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n755), .B2(new_n376), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n361), .B1(new_n202), .B2(new_n763), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n758), .C1(new_n781), .C2(new_n768), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n929), .A2(new_n762), .B1(new_n271), .B2(new_n745), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n832), .B(new_n1122), .C1(G107), .C2(new_n749), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n364), .B1(new_n742), .B2(new_n492), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G294), .B2(new_n759), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n770), .A3(new_n1040), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n787), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n373), .B2(new_n835), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n790), .B(new_n1128), .C1(new_n1084), .C2(new_n801), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT110), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1082), .B1(new_n1100), .B2(new_n1083), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n950), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1107), .A2(new_n1131), .A3(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(new_n881), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n890), .C2(new_n1085), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT115), .B1(new_n619), .B2(new_n392), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n403), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n381), .A2(new_n856), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n403), .A2(new_n1140), .ZN(new_n1147));
  AOI211_X1 g0947(.A(KEYINPUT115), .B(new_n392), .C1(new_n400), .C2(new_n402), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n908), .B2(G330), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n907), .A2(new_n905), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n906), .A2(new_n903), .A3(new_n895), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n1150), .A3(G330), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1138), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(G330), .A3(new_n1153), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1150), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n892), .A3(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n950), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n835), .A2(new_n202), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n749), .A2(G132), .B1(new_n817), .B2(G137), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT113), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n929), .A2(new_n1120), .B1(new_n755), .B2(new_n1110), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G150), .B2(new_n779), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n1108), .C2(new_n742), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT114), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G33), .B1(new_n759), .B2(G124), .ZN(new_n1172));
  AOI21_X1  g0972(.A(G41), .B1(new_n773), .B2(G159), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n202), .B1(new_n261), .B2(G41), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n763), .A2(new_n207), .B1(new_n762), .B2(new_n758), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1177), .A2(new_n275), .A3(new_n1042), .A4(new_n1012), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT111), .Z(new_n1179));
  AOI22_X1  g0979(.A1(new_n775), .A2(G107), .B1(new_n749), .B2(G97), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n492), .B2(new_n929), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G68), .B2(new_n779), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n343), .C2(new_n745), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT112), .B(KEYINPUT58), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1174), .A2(new_n1175), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n791), .B1(new_n1186), .B2(new_n788), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1163), .B(new_n1187), .C1(new_n1150), .C2(new_n801), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1106), .A2(new_n1072), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n1161), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1021), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1161), .A3(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G375));
  NAND3_X1  g0996(.A1(new_n1070), .A2(KEYINPUT116), .A3(new_n950), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT116), .B1(new_n1070), .B2(new_n950), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n929), .A2(new_n1112), .B1(new_n924), .B2(new_n742), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n477), .B1(new_n763), .B2(new_n207), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n755), .A2(new_n781), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1108), .B2(new_n758), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1201), .B(new_n1205), .C1(new_n749), .C2(new_n1109), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n202), .B2(new_n768), .C1(new_n376), .C2(new_n745), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n929), .A2(new_n764), .B1(new_n214), .B2(new_n745), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G116), .B2(new_n749), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1009), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n361), .B1(new_n775), .B2(G283), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n756), .A2(G97), .B1(new_n773), .B2(G77), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n758), .A2(new_n938), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(new_n788), .B1(new_n222), .B2(new_n835), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n790), .B(new_n1216), .C1(new_n855), .C2(new_n801), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1061), .A2(new_n1071), .A3(new_n1069), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1073), .A2(new_n971), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1200), .A2(new_n1217), .A3(new_n1219), .ZN(G381));
  NOR3_X1   g1020(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(G407));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1223), .B2(new_n671), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G407), .A2(new_n1226), .ZN(G409));
  AOI22_X1  g1027(.A1(new_n1072), .A2(new_n1106), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n971), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G378), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1022), .B1(new_n1228), .B2(KEYINPUT57), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1194), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1230), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT117), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1159), .A2(new_n892), .A3(new_n1154), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n892), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1071), .B1(new_n1133), .B2(new_n1070), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1192), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1022), .A3(new_n1194), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(KEYINPUT117), .A3(G378), .A4(new_n1230), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1231), .B1(new_n1236), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G384), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1218), .A2(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1061), .A2(new_n1071), .A3(new_n1069), .A4(KEYINPUT60), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1073), .A3(new_n1022), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1070), .A2(new_n950), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT116), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1217), .A3(new_n1197), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1245), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1200), .A2(new_n1249), .A3(G384), .A4(new_n1217), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1255), .A2(KEYINPUT118), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT118), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1225), .A2(G343), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1244), .A2(new_n1260), .A3(KEYINPUT62), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1231), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT117), .B1(new_n1195), .B2(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1243), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1261), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT124), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1244), .A2(new_n1269), .A3(new_n1261), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1259), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1262), .B1(new_n1271), .B2(KEYINPUT62), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1266), .A2(KEYINPUT124), .A3(new_n1267), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1269), .B1(new_n1244), .B2(new_n1261), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1261), .A2(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT119), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1278), .B1(new_n1281), .B2(KEYINPUT119), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1274), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1283), .A2(KEYINPUT125), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1272), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1288));
  XOR2_X1   g1088(.A(G393), .B(G396), .Z(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(KEYINPUT120), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT121), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  OR3_X1    g1094(.A1(G387), .A2(new_n1294), .A3(KEYINPUT122), .ZN(new_n1295));
  AND2_X1   g1095(.A1(G387), .A2(new_n1294), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT122), .B1(G387), .B2(new_n1294), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1293), .B(new_n1295), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  AND3_X1   g1098(.A1(G387), .A2(KEYINPUT123), .A3(G390), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G390), .B1(G387), .B2(KEYINPUT123), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1290), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1292), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1272), .B(new_n1304), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1288), .A2(new_n1303), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1260), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1307), .B2(KEYINPUT63), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1244), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1282), .B1(new_n1261), .B2(new_n1244), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1310), .A2(KEYINPUT63), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1308), .B(new_n1302), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(new_n1312), .ZN(G405));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  INV_X1    g1114(.A(G378), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1236), .A2(new_n1243), .B1(new_n1315), .B2(G375), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1275), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1260), .B2(new_n1316), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1302), .A2(new_n1314), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1302), .A2(new_n1318), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1314), .B1(new_n1302), .B2(new_n1318), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(G402));
endmodule


