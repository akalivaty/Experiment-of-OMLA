

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X2 U321 ( .A(KEYINPUT37), .B(n494), .ZN(n519) );
  XNOR2_X1 U322 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U323 ( .A(n310), .B(n410), .Z(n535) );
  NOR2_X1 U324 ( .A1(n382), .A2(n575), .ZN(n399) );
  XNOR2_X1 U325 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U326 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n426) );
  XNOR2_X1 U327 ( .A(n330), .B(G29GAT), .ZN(n331) );
  XNOR2_X1 U328 ( .A(n427), .B(n426), .ZN(n449) );
  XNOR2_X1 U329 ( .A(n332), .B(n331), .ZN(n334) );
  NOR2_X1 U330 ( .A1(n535), .A2(n451), .ZN(n569) );
  XOR2_X1 U331 ( .A(n448), .B(n447), .Z(n520) );
  XNOR2_X1 U332 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n290) );
  XNOR2_X1 U335 ( .A(G15GAT), .B(KEYINPUT92), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U337 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n292) );
  XNOR2_X1 U338 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U340 ( .A(n294), .B(n293), .Z(n306) );
  XNOR2_X1 U341 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n295), .B(KEYINPUT86), .ZN(n296) );
  XOR2_X1 U343 ( .A(n296), .B(G134GAT), .Z(n298) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n297) );
  XOR2_X1 U345 ( .A(n298), .B(n297), .Z(n446) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n368) );
  XOR2_X1 U347 ( .A(G176GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G43GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U350 ( .A(n368), .B(n301), .Z(n303) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U352 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U353 ( .A(n446), .B(n304), .Z(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U355 ( .A(G183GAT), .B(G190GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(KEYINPUT19), .B(n309), .Z(n410) );
  XOR2_X1 U359 ( .A(KEYINPUT3), .B(KEYINPUT93), .Z(n312) );
  XNOR2_X1 U360 ( .A(G162GAT), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U362 ( .A(KEYINPUT2), .B(n313), .Z(n428) );
  XOR2_X1 U363 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n315) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G197GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n428), .B(n316), .ZN(n327) );
  XOR2_X1 U367 ( .A(KEYINPUT21), .B(G211GAT), .Z(n318) );
  XNOR2_X1 U368 ( .A(G204GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n415) );
  XOR2_X1 U370 ( .A(G141GAT), .B(G22GAT), .Z(n386) );
  XOR2_X1 U371 ( .A(n415), .B(n386), .Z(n320) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U374 ( .A(n321), .B(KEYINPUT24), .Z(n325) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n377) );
  XNOR2_X1 U378 ( .A(n377), .B(KEYINPUT94), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n474) );
  XOR2_X1 U381 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n329) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n347) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n332) );
  INV_X1 U385 ( .A(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U386 ( .A(G43GAT), .B(G50GAT), .ZN(n333) );
  XOR2_X1 U387 ( .A(n334), .B(n333), .Z(n397) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(KEYINPUT76), .ZN(n369) );
  XOR2_X1 U390 ( .A(n397), .B(n369), .Z(n343) );
  XOR2_X1 U391 ( .A(KEYINPUT67), .B(KEYINPUT79), .Z(n337) );
  XNOR2_X1 U392 ( .A(G134GAT), .B(G162GAT), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n339) );
  XOR2_X1 U394 ( .A(G190GAT), .B(G218GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n340) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n558) );
  XNOR2_X1 U400 ( .A(n558), .B(KEYINPUT36), .ZN(n491) );
  XOR2_X1 U401 ( .A(KEYINPUT82), .B(G64GAT), .Z(n349) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U404 ( .A(n350), .B(G71GAT), .Z(n352) );
  XOR2_X1 U405 ( .A(G15GAT), .B(G1GAT), .Z(n385) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(n385), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(G211GAT), .Z(n354) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n356) );
  XNOR2_X1 U412 ( .A(G127GAT), .B(G155GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U415 ( .A(KEYINPUT13), .B(G57GAT), .Z(n367) );
  XOR2_X1 U416 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n360) );
  XNOR2_X1 U417 ( .A(G183GAT), .B(KEYINPUT81), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n367), .B(n361), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n580) );
  INV_X1 U422 ( .A(n580), .ZN(n554) );
  NOR2_X1 U423 ( .A1(n491), .A2(n554), .ZN(n366) );
  XOR2_X1 U424 ( .A(n366), .B(KEYINPUT45), .Z(n382) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U426 ( .A(n369), .B(G204GAT), .Z(n371) );
  NAND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U429 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT31), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U433 ( .A(G176GAT), .B(G92GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n376), .B(G64GAT), .ZN(n418) );
  XNOR2_X1 U435 ( .A(n377), .B(n418), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n575) );
  XOR2_X1 U438 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n384) );
  XNOR2_X1 U439 ( .A(KEYINPUT73), .B(G113GAT), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U441 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n388) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U445 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U447 ( .A(n393), .B(KEYINPUT70), .Z(n396) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(G8GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(G197GAT), .ZN(n420) );
  XNOR2_X1 U450 ( .A(n420), .B(KEYINPUT30), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U452 ( .A(n398), .B(n397), .Z(n548) );
  INV_X1 U453 ( .A(n548), .ZN(n571) );
  XOR2_X1 U454 ( .A(KEYINPUT74), .B(n571), .Z(n536) );
  NAND2_X1 U455 ( .A1(n399), .A2(n536), .ZN(n407) );
  INV_X1 U456 ( .A(n558), .ZN(n542) );
  XOR2_X1 U457 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n402) );
  XNOR2_X1 U458 ( .A(n575), .B(KEYINPUT65), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n400), .B(KEYINPUT41), .ZN(n566) );
  NAND2_X1 U460 ( .A1(n566), .A2(n571), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n403), .A2(n554), .ZN(n404) );
  NOR2_X1 U463 ( .A1(n542), .A2(n404), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n405), .B(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U465 ( .A1(n407), .A2(n406), .ZN(n409) );
  XNOR2_X1 U466 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n530) );
  INV_X1 U468 ( .A(n410), .ZN(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n412) );
  XNOR2_X1 U470 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U472 ( .A(n414), .B(n413), .Z(n424) );
  XOR2_X1 U473 ( .A(n415), .B(KEYINPUT80), .Z(n417) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U476 ( .A(n419), .B(n418), .Z(n422) );
  XNOR2_X1 U477 ( .A(G36GAT), .B(n420), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n522) );
  INV_X1 U480 ( .A(n522), .ZN(n425) );
  NAND2_X1 U481 ( .A1(n530), .A2(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT99), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(KEYINPUT98), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n431), .B(KEYINPUT6), .Z(n439) );
  XOR2_X1 U486 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n433) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U489 ( .A(G148GAT), .B(G57GAT), .Z(n435) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n441) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(G85GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n448) );
  INV_X1 U500 ( .A(n446), .ZN(n447) );
  NAND2_X1 U501 ( .A1(n449), .A2(n520), .ZN(n457) );
  NOR2_X1 U502 ( .A1(n474), .A2(n457), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U504 ( .A1(n569), .A2(n542), .ZN(n453) );
  INV_X1 U505 ( .A(G218GAT), .ZN(n462) );
  XOR2_X1 U506 ( .A(KEYINPUT106), .B(KEYINPUT26), .Z(n455) );
  NAND2_X1 U507 ( .A1(n474), .A2(n535), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n547) );
  INV_X1 U509 ( .A(n547), .ZN(n456) );
  NOR2_X1 U510 ( .A1(n457), .A2(n456), .ZN(n581) );
  INV_X1 U511 ( .A(n581), .ZN(n458) );
  NOR2_X1 U512 ( .A1(n491), .A2(n458), .ZN(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(G1355GAT) );
  XOR2_X1 U516 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n464) );
  NAND2_X1 U517 ( .A1(n580), .A2(n558), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n464), .B(n463), .ZN(n480) );
  NOR2_X1 U519 ( .A1(n535), .A2(n522), .ZN(n465) );
  NOR2_X1 U520 ( .A1(n474), .A2(n465), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT25), .ZN(n468) );
  XOR2_X1 U522 ( .A(n522), .B(KEYINPUT27), .Z(n471) );
  NAND2_X1 U523 ( .A1(n547), .A2(n471), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n520), .A2(n469), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT107), .B(n470), .Z(n479) );
  INV_X1 U527 ( .A(n471), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n472), .A2(n520), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT104), .ZN(n531) );
  XOR2_X1 U530 ( .A(n474), .B(KEYINPUT68), .Z(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT28), .B(n475), .ZN(n533) );
  NAND2_X1 U532 ( .A1(n531), .A2(n533), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT105), .B(n476), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n535), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n493) );
  AND2_X1 U536 ( .A1(n480), .A2(n493), .ZN(n509) );
  NOR2_X1 U537 ( .A1(n575), .A2(n536), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n481), .B(KEYINPUT78), .ZN(n495) );
  NAND2_X1 U539 ( .A1(n509), .A2(n495), .ZN(n489) );
  NOR2_X1 U540 ( .A1(n520), .A2(n489), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT108), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U543 ( .A(G1GAT), .B(n484), .Z(G1324GAT) );
  NOR2_X1 U544 ( .A1(n522), .A2(n489), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT109), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1325GAT) );
  NOR2_X1 U547 ( .A1(n535), .A2(n489), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n533), .A2(n489), .ZN(n490) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U552 ( .A1(n491), .A2(n580), .ZN(n492) );
  NAND2_X1 U553 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n519), .A2(n495), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(KEYINPUT110), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n502) );
  NOR2_X1 U557 ( .A1(n520), .A2(n502), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  BUF_X1 U560 ( .A(n502), .Z(n506) );
  NOR2_X1 U561 ( .A1(n522), .A2(n506), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(KEYINPUT111), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n535), .A2(n502), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U567 ( .A(G43GAT), .B(n505), .Z(G1330GAT) );
  NOR2_X1 U568 ( .A1(n533), .A2(n506), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT113), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  INV_X1 U571 ( .A(n566), .ZN(n550) );
  NOR2_X1 U572 ( .A1(n571), .A2(n550), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n518), .A2(n509), .ZN(n515) );
  NOR2_X1 U574 ( .A1(n520), .A2(n515), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n522), .A2(n515), .ZN(n512) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n535), .A2(n515), .ZN(n513) );
  XOR2_X1 U580 ( .A(KEYINPUT114), .B(n513), .Z(n514) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U582 ( .A1(n533), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n520), .A2(n526), .ZN(n521) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n535), .A2(n526), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n533), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(n532), .Z(n546) );
  NAND2_X1 U599 ( .A1(n533), .A2(n546), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n543) );
  INV_X1 U601 ( .A(n536), .ZN(n561) );
  NAND2_X1 U602 ( .A1(n543), .A2(n561), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U605 ( .A1(n543), .A2(n566), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n543), .A2(n580), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n548), .A2(n557), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n557), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n557), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n559), .Z(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n569), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .Z(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n580), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n573) );
  NAND2_X1 U637 ( .A1(n581), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n579) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT124), .Z(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
endmodule

