//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G120gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT1), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G127gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G134gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n222), .A3(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n217), .A2(new_n222), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n225), .B1(new_n230), .B2(new_n215), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n217), .A2(new_n222), .A3(new_n228), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n217), .B2(new_n222), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n225), .B(new_n215), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G141gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G148gat), .ZN(new_n238));
  INV_X1    g037(.A(G148gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G141gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n238), .A2(new_n240), .B1(KEYINPUT2), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G155gat), .B(G162gat), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(KEYINPUT2), .ZN(new_n246));
  AND4_X1   g045(.A1(KEYINPUT72), .A2(new_n245), .A3(new_n243), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT72), .B1(new_n242), .B2(new_n243), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n210), .B1(new_n236), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n223), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n251), .A2(new_n215), .A3(new_n219), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n215), .B1(new_n232), .B2(new_n233), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n242), .A2(new_n243), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n245), .A2(new_n243), .A3(new_n246), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n242), .A2(KEYINPUT72), .A3(new_n243), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n255), .A2(KEYINPUT75), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n231), .A2(new_n235), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n224), .B(new_n244), .C1(new_n248), .C2(new_n247), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT74), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n234), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n252), .A2(new_n256), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n209), .B1(new_n263), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n244), .C1(new_n247), .C2(new_n248), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n236), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n277), .A2(new_n208), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT4), .B1(new_n266), .B2(new_n271), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n264), .A2(new_n265), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n278), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n283), .A3(KEYINPUT5), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n208), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n271), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n280), .A2(new_n281), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n290), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(KEYINPUT6), .B(new_n207), .C1(new_n285), .C2(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n290), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT76), .B1(new_n289), .B2(new_n290), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n287), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n284), .A3(new_n206), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n206), .B1(new_n299), .B2(new_n284), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n305));
  INV_X1    g104(.A(KEYINPUT37), .ZN(new_n306));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(G183gat), .A3(G190gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G183gat), .B(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n309), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n308), .B1(new_n312), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n314), .A2(KEYINPUT65), .A3(new_n315), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT65), .B1(new_n314), .B2(new_n315), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(KEYINPUT64), .A2(new_n319), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n310), .ZN(new_n326));
  XOR2_X1   g125(.A(G183gat), .B(G190gat), .Z(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(KEYINPUT24), .ZN(new_n328));
  INV_X1    g127(.A(new_n318), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT25), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n335), .B(KEYINPUT28), .Z(new_n336));
  INV_X1    g135(.A(new_n313), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT26), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n315), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n313), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n325), .A2(new_n332), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n307), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n341), .ZN(new_n344));
  INV_X1    g143(.A(new_n323), .ZN(new_n345));
  INV_X1    g144(.A(new_n320), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n314), .A2(KEYINPUT65), .A3(new_n315), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n330), .B2(new_n331), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n319), .A2(KEYINPUT64), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n307), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G197gat), .A2(G204gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n361), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n306), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n342), .A2(KEYINPUT70), .A3(new_n307), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n351), .B2(new_n352), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n369), .B(new_n343), .C1(new_n370), .C2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n305), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n367), .B(new_n343), .C1(new_n370), .C2(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n352), .B1(new_n351), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n342), .A2(new_n307), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n369), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n383), .A3(new_n377), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n202), .B1(new_n304), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n385), .A2(new_n378), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n367), .B1(new_n343), .B2(new_n353), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n353), .A2(KEYINPUT70), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n351), .A2(new_n371), .A3(new_n352), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n381), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n394), .B2(new_n367), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n390), .A2(new_n374), .B1(new_n395), .B2(new_n377), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n207), .B1(new_n285), .B2(new_n295), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n301), .A3(new_n300), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT84), .A4(new_n296), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n390), .B1(new_n306), .B2(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n305), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n389), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT39), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n263), .A2(new_n272), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n208), .ZN(new_n405));
  INV_X1    g204(.A(new_n277), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n293), .B2(new_n294), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n208), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n277), .B1(new_n297), .B2(new_n298), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n403), .A3(new_n209), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n408), .A2(KEYINPUT40), .A3(new_n206), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n379), .A2(new_n383), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n378), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n383), .A4(new_n377), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n408), .A2(new_n206), .A3(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT40), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n303), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(KEYINPUT78), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n367), .A2(new_n380), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n275), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n249), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n367), .B1(new_n276), .B2(new_n380), .ZN(new_n432));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT29), .B1(new_n261), .B2(new_n275), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT3), .B1(new_n367), .B2(new_n380), .ZN(new_n437));
  OAI22_X1  g236(.A1(new_n436), .A2(new_n367), .B1(new_n261), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT80), .B1(new_n438), .B2(new_n433), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n437), .A2(new_n261), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT80), .B(new_n433), .C1(new_n432), .C2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n435), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G22gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n433), .B1(new_n432), .B2(new_n440), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(G22gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n435), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n426), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT79), .B(new_n425), .C1(new_n444), .C2(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n423), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI221_X4 g254(.A(G22gat), .B1(new_n431), .B2(new_n434), .C1(new_n447), .C2(new_n441), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n448), .B2(new_n435), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n425), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n452), .A3(new_n426), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n422), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n418), .A2(new_n421), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n402), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n301), .B(new_n300), .C1(new_n303), .C2(new_n464), .ZN(new_n465));
  AOI211_X1 g264(.A(KEYINPUT77), .B(new_n206), .C1(new_n299), .C2(new_n284), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n296), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n415), .A2(new_n468), .A3(new_n416), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n413), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n415), .B2(new_n416), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n459), .A2(new_n422), .A3(new_n460), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n422), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n342), .A2(new_n236), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n351), .A2(new_n255), .ZN(new_n478));
  INV_X1    g277(.A(G227gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G15gat), .B(G43gat), .Z(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n488), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n482), .B(KEYINPUT32), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n478), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n479), .B2(new_n480), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT34), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n493), .B(new_n496), .C1(new_n479), .C2(new_n480), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n489), .A2(new_n495), .A3(new_n497), .A4(new_n491), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT36), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n492), .A2(new_n498), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n473), .A2(new_n476), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n463), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n500), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n476), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(KEYINPUT35), .A3(new_n467), .A4(new_n472), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n455), .A2(new_n461), .B1(new_n502), .B2(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(new_n417), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n304), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n304), .A2(KEYINPUT85), .A3(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n508), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT86), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n526), .A2(KEYINPUT14), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n524), .B2(new_n525), .ZN(new_n530));
  NAND3_X1  g329(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(KEYINPUT14), .C2(new_n527), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  XOR2_X1   g332(.A(G43gat), .B(G50gat), .Z(new_n534));
  AOI211_X1 g333(.A(new_n528), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n534), .A2(new_n533), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT16), .A3(new_n543), .ZN(new_n544));
  OAI221_X1 g343(.A(new_n544), .B1(KEYINPUT89), .B2(G8gat), .C1(new_n543), .C2(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n539), .B(KEYINPUT88), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT17), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n537), .A2(KEYINPUT17), .A3(new_n538), .ZN(new_n551));
  INV_X1    g350(.A(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n522), .B(new_n548), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n541), .B(new_n552), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n522), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G197gat), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT11), .B(G169gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT12), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n556), .A2(new_n569), .A3(new_n560), .A4(new_n561), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n521), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(KEYINPUT8), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G99gat), .B(G106gat), .Z(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT93), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n551), .B(new_n589), .C1(new_n549), .C2(KEYINPUT17), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n541), .A2(new_n591), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(new_n595), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n576), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT94), .B(new_n576), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(new_n576), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n594), .B2(new_n596), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT9), .ZN(new_n609));
  INV_X1    g408(.A(G57gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G64gat), .ZN(new_n611));
  INV_X1    g410(.A(G64gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G57gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n615));
  INV_X1    g414(.A(G71gat), .ZN(new_n616));
  INV_X1    g415(.A(G78gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n618), .B2(new_n609), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n611), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n615), .B1(new_n614), .B2(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G127gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n552), .B1(new_n629), .B2(new_n628), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  INV_X1    g435(.A(G155gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G183gat), .B(G211gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n635), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n589), .A2(new_n643), .A3(new_n628), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n589), .A2(new_n628), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n585), .A2(new_n587), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(new_n628), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n645), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT96), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n644), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G230gat), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n480), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n642), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n644), .ZN(new_n657));
  INV_X1    g456(.A(new_n652), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n648), .A2(new_n651), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n655), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(KEYINPUT97), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n661), .B1(new_n645), .B2(new_n647), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  NOR2_X1   g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n656), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n655), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n671), .B2(new_n663), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n608), .A2(new_n641), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n572), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n467), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n543), .ZN(G1324gat));
  INV_X1    g476(.A(G8gat), .ZN(new_n678));
  INV_X1    g477(.A(new_n675), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n417), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n678), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n675), .A2(new_n513), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n502), .A2(new_n505), .ZN(new_n686));
  AOI21_X1  g485(.A(G15gat), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n506), .A2(new_n501), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT101), .Z(new_n691));
  AOI21_X1  g490(.A(new_n687), .B1(new_n679), .B2(new_n691), .ZN(G1326gat));
  AND2_X1   g491(.A1(new_n572), .A2(new_n476), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n674), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT102), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n608), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n508), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n463), .A2(new_n507), .A3(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n511), .A2(new_n520), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n699), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n521), .B2(new_n608), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n673), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n641), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n568), .A2(new_n570), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT103), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n467), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n521), .A2(new_n608), .A3(new_n713), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(G29gat), .A3(new_n467), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT45), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1328gat));
  OAI21_X1  g519(.A(G36gat), .B1(new_n715), .B2(new_n513), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n717), .A2(G36gat), .A3(new_n513), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1329gat));
  NAND2_X1  g523(.A1(new_n689), .A2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n686), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n715), .A2(new_n725), .B1(G43gat), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g528(.A(new_n476), .ZN(new_n730));
  OAI21_X1  g529(.A(G50gat), .B1(new_n715), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n608), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n711), .A2(new_n732), .A3(G50gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n693), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT48), .Z(G1331gat));
  AOI21_X1  g535(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  INV_X1    g537(.A(new_n641), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n732), .A2(new_n712), .A3(new_n739), .A4(new_n673), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n738), .B1(new_n737), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n467), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(new_n610), .ZN(G1332gat));
  INV_X1    g544(.A(new_n743), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT49), .B(G64gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n417), .A3(new_n747), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n743), .A2(new_n513), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n746), .A2(KEYINPUT107), .A3(new_n686), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n743), .B2(new_n726), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n616), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n746), .A2(G71gat), .A3(new_n689), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n754), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1334gat));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n730), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(new_n617), .ZN(G1335gat));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n571), .B2(new_n739), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n568), .A2(KEYINPUT109), .A3(new_n570), .A4(new_n641), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n765), .B2(new_n673), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n767), .B(new_n710), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n709), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n467), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n608), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n737), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n467), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n673), .A2(new_n580), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n771), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT111), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n770), .B2(new_n513), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT113), .B1(new_n737), .B2(new_n772), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n774), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n737), .C2(new_n772), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n710), .A2(G92gat), .A3(new_n513), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT112), .Z(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n775), .B2(new_n785), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n781), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n770), .B2(new_n688), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n710), .A2(G99gat), .A3(new_n726), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n776), .B2(new_n797), .ZN(G1338gat));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n673), .A2(new_n799), .A3(new_n476), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n775), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n476), .B(new_n769), .C1(new_n706), .C2(new_n708), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n801), .B(KEYINPUT116), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n783), .A2(new_n807), .A3(new_n784), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n805), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT117), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n811), .B(new_n803), .C1(new_n808), .C2(new_n805), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n806), .B(KEYINPUT118), .C1(new_n810), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(new_n668), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n671), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n655), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT119), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n656), .A2(KEYINPUT54), .A3(new_n662), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n820), .B(KEYINPUT55), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n826), .A2(new_n571), .A3(new_n670), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n557), .A2(new_n559), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n548), .B1(new_n550), .B2(new_n553), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(G229gat), .A3(G233gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n829), .A2(new_n830), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n566), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n570), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n673), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n608), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n837), .A2(new_n608), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n827), .A2(new_n670), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(new_n826), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n641), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n674), .A2(new_n712), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(new_n777), .A3(new_n510), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n513), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n571), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n512), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n777), .A2(new_n513), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n712), .A2(new_n213), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(G1340gat));
  AOI21_X1  g652(.A(G120gat), .B1(new_n847), .B2(new_n673), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n710), .A2(new_n211), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n851), .B2(new_n855), .ZN(G1341gat));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n221), .A3(new_n739), .ZN(new_n857));
  INV_X1    g656(.A(new_n851), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n858), .B2(new_n641), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1342gat));
  NAND4_X1  g659(.A1(new_n846), .A2(new_n216), .A3(new_n513), .A4(new_n608), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n858), .B2(new_n732), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NOR2_X1   g664(.A1(new_n689), .A2(new_n850), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT121), .Z(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n730), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n844), .B1(new_n843), .B2(KEYINPUT122), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n840), .A2(new_n841), .A3(new_n826), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n712), .B1(new_n825), .B2(new_n824), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n873), .A2(new_n841), .B1(new_n673), .B2(new_n837), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(new_n608), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n871), .B1(new_n875), .B2(new_n641), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n869), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n875), .A2(new_n641), .B1(new_n712), .B2(new_n674), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n868), .B1(new_n878), .B2(new_n730), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n867), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n237), .B1(new_n880), .B2(new_n571), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n689), .A2(new_n730), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n845), .A2(new_n777), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n417), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n237), .A3(new_n571), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT58), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n712), .B(new_n867), .C1(new_n877), .C2(new_n879), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n885), .B(new_n888), .C1(new_n889), .C2(new_n237), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n239), .A3(new_n673), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n239), .C1(new_n880), .C2(new_n673), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n867), .A2(new_n710), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n845), .A2(new_n476), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n868), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n845), .B2(new_n476), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n892), .B1(new_n893), .B2(new_n900), .ZN(G1345gat));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n637), .A3(new_n739), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n880), .A2(new_n739), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n637), .ZN(G1346gat));
  OR4_X1    g703(.A1(G162gat), .A2(new_n883), .A3(new_n417), .A4(new_n732), .ZN(new_n905));
  AOI211_X1 g704(.A(new_n732), .B(new_n867), .C1(new_n877), .C2(new_n879), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  OAI21_X1  g706(.A(G162gat), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n880), .A2(new_n907), .A3(new_n608), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n777), .A2(new_n513), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n845), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n510), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n571), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n911), .B(KEYINPUT124), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n849), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n571), .A2(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  INV_X1    g717(.A(new_n916), .ZN(new_n919));
  OAI21_X1  g718(.A(G176gat), .B1(new_n919), .B2(new_n710), .ZN(new_n920));
  INV_X1    g719(.A(G176gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n921), .A3(new_n673), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(G183gat), .B1(new_n919), .B2(new_n641), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n913), .A2(new_n333), .A3(new_n739), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n334), .A3(new_n608), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n608), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(G190gat), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT61), .B(new_n334), .C1(new_n916), .C2(new_n608), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n712), .A2(G197gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n912), .A2(new_n882), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT126), .Z(new_n938));
  NOR2_X1   g737(.A1(new_n915), .A2(new_n689), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n897), .B2(new_n898), .ZN(new_n940));
  OAI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n712), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(new_n941), .ZN(G1352gat));
  OAI21_X1  g741(.A(G204gat), .B1(new_n940), .B2(new_n710), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n710), .A2(G204gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n912), .A2(new_n882), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n912), .A2(new_n948), .A3(new_n882), .A4(new_n944), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n946), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(G1353gat));
  AND2_X1   g751(.A1(new_n912), .A2(new_n882), .ZN(new_n953));
  INV_X1    g752(.A(G211gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(new_n739), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n739), .B(new_n939), .C1(new_n897), .C2(new_n898), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n940), .B2(new_n732), .ZN(new_n960));
  INV_X1    g759(.A(G218gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n961), .A3(new_n608), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1355gat));
endmodule


