//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT23), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(new_n201), .C1(new_n197), .C2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G110), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  XNOR2_X1  g019(.A(G119), .B(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT74), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT16), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n213), .A2(KEYINPUT16), .A3(G140), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n213), .A2(KEYINPUT16), .A3(G140), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT74), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n209), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n219), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n222), .B2(KEYINPUT16), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(G146), .C1(new_n223), .C2(new_n210), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n208), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI22_X1  g039(.A1(new_n203), .A2(G110), .B1(new_n206), .B2(new_n205), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n209), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n226), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n195), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n224), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n207), .A3(new_n204), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n224), .A3(new_n227), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n194), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n233), .A3(new_n188), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n229), .A2(new_n233), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n190), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n189), .A2(G902), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n229), .A2(new_n233), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g057(.A(G116), .B(G119), .Z(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT30), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n209), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G143), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G146), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n250), .B2(G146), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n251), .A2(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G137), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .A3(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(G137), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT67), .B(G131), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n265), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G131), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT68), .B1(new_n259), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n276), .A3(G146), .ZN(new_n277));
  INV_X1    g091(.A(new_n253), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n276), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n248), .B1(new_n280), .B2(new_n209), .ZN(new_n281));
  INV_X1    g095(.A(new_n255), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n266), .A2(new_n267), .B1(G131), .B2(new_n270), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n273), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G131), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n268), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n278), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT0), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n257), .A3(KEYINPUT64), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(KEYINPUT0), .B2(G128), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n296), .A2(new_n298), .B1(KEYINPUT0), .B2(G128), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n251), .A2(KEYINPUT66), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT66), .B1(new_n251), .B2(new_n299), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n290), .B(new_n294), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n247), .B1(new_n287), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n283), .A2(new_n284), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n247), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n246), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n246), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n285), .B1(new_n283), .B2(new_n284), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n302), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT69), .B(G237), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(new_n192), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G210), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n316), .A3(G210), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT26), .B(G101), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT70), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n311), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n307), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n307), .A2(new_n323), .A3(KEYINPUT31), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n302), .A2(new_n304), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT71), .A3(new_n246), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n311), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT71), .B1(new_n331), .B2(new_n246), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT28), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n331), .B2(new_n246), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n321), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(G902), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G472), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT32), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n328), .A2(new_n329), .B1(new_n338), .B2(new_n339), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n345));
  NOR4_X1   g159(.A1(new_n344), .A2(new_n345), .A3(G472), .A4(G902), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n308), .B1(new_n349), .B2(new_n305), .ZN(new_n350));
  INV_X1    g164(.A(new_n311), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT72), .B1(new_n352), .B2(new_n321), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n335), .A2(new_n337), .A3(new_n321), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n339), .C1(new_n350), .C2(new_n351), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n246), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n311), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT28), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(new_n337), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n339), .A2(new_n354), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G472), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n243), .B1(new_n347), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n297), .A2(KEYINPUT0), .A3(G128), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT64), .B1(new_n295), .B2(new_n257), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n292), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n281), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n251), .A2(KEYINPUT66), .A3(new_n299), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(G101), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n376), .A2(new_n379), .A3(new_n385), .A4(new_n380), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n374), .A2(new_n294), .A3(new_n383), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n277), .A2(new_n278), .A3(new_n258), .ZN(new_n390));
  AOI21_X1  g204(.A(G146), .B1(new_n274), .B2(new_n276), .ZN(new_n391));
  OAI21_X1  g205(.A(G128), .B1(new_n391), .B2(new_n254), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n291), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT76), .B1(new_n375), .B2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n380), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n375), .A2(KEYINPUT76), .A3(G107), .ZN(new_n396));
  OAI21_X1  g210(.A(G101), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n386), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n389), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n290), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n251), .A2(new_n255), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n389), .B1(new_n401), .B2(new_n279), .ZN(new_n402));
  INV_X1    g216(.A(new_n398), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n388), .A2(new_n399), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n387), .A2(new_n383), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n293), .B1(new_n372), .B2(new_n373), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n408), .A2(new_n409), .B1(new_n403), .B2(new_n402), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(KEYINPUT77), .A3(new_n400), .A4(new_n399), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n290), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT75), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n192), .A2(G227), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n393), .A2(new_n398), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n403), .A2(new_n283), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n290), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT12), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n419), .B1(new_n407), .B2(new_n411), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI211_X1 g242(.A(KEYINPUT78), .B(new_n419), .C1(new_n407), .C2(new_n411), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n420), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G469), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n188), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n412), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n419), .B1(new_n414), .B2(new_n426), .ZN(new_n434));
  OAI21_X1  g248(.A(G469), .B1(new_n434), .B2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G221), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n439), .B2(new_n188), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT79), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n246), .A2(new_n387), .A3(new_n383), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n244), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G116), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n456), .A2(KEYINPUT5), .A3(G119), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n455), .A2(G113), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n244), .A2(new_n245), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n403), .A3(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n246), .A2(new_n387), .A3(KEYINPUT80), .A4(new_n383), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n453), .A2(new_n465), .A3(new_n462), .A4(new_n463), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n259), .A2(new_n213), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n409), .B2(new_n213), .ZN(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n475), .A3(new_n466), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n403), .B1(new_n461), .B2(new_n460), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n465), .B(KEYINPUT8), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n478), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n409), .A2(new_n213), .ZN(new_n484));
  INV_X1    g298(.A(new_n473), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(KEYINPUT7), .A3(new_n485), .A4(new_n470), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n473), .B1(KEYINPUT83), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(KEYINPUT83), .B2(new_n487), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n471), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n483), .A2(new_n486), .A3(new_n468), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n188), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n450), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(new_n188), .A3(new_n449), .A4(new_n491), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n448), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(G113), .B(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(new_n375), .ZN(new_n498));
  AND2_X1   g312(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n499));
  NOR2_X1   g313(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n222), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n222), .B2(new_n500), .ZN(new_n502));
  AND2_X1   g316(.A1(KEYINPUT69), .A2(G237), .ZN(new_n503));
  NOR2_X1   g317(.A1(KEYINPUT69), .A2(G237), .ZN(new_n504));
  OAI211_X1 g318(.A(G214), .B(new_n192), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n274), .A2(new_n276), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(G143), .B1(new_n275), .B2(KEYINPUT84), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n312), .A2(G214), .A3(new_n192), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n267), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  OAI221_X1 g327(.A(new_n224), .B1(G146), .B2(new_n502), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n510), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n222), .B(new_n209), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT18), .A4(G131), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n498), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n512), .A2(new_n513), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n523), .A2(new_n524), .B1(new_n230), .B2(KEYINPUT86), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n220), .A2(new_n224), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n521), .B1(new_n530), .B2(new_n498), .ZN(new_n531));
  NOR2_X1   g345(.A1(G475), .A2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT20), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n230), .A2(KEYINPUT86), .ZN(new_n535));
  INV_X1    g349(.A(new_n513), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n524), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n535), .A2(new_n538), .A3(new_n527), .A4(new_n528), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n498), .A3(new_n520), .ZN(new_n540));
  INV_X1    g354(.A(new_n521), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n532), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n539), .A2(new_n498), .A3(new_n520), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n498), .B1(new_n539), .B2(new_n520), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n188), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n534), .A2(new_n544), .B1(G475), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT87), .ZN(new_n549));
  INV_X1    g363(.A(G122), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(G116), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n456), .A2(KEYINPUT87), .A3(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(G116), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(KEYINPUT14), .ZN(new_n557));
  OAI21_X1  g371(.A(G107), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n257), .A2(G143), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n280), .B2(new_n257), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G134), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n261), .B(new_n559), .C1(new_n280), .C2(new_n257), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n378), .A3(new_n555), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n558), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n555), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G107), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n250), .A2(new_n569), .A3(G128), .ZN(new_n570));
  OAI211_X1 g384(.A(G134), .B(new_n570), .C1(new_n560), .C2(new_n569), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n571), .A3(new_n562), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n438), .A2(new_n187), .A3(G953), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n565), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n565), .A2(new_n572), .ZN(new_n578));
  INV_X1    g392(.A(new_n573), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n188), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n581), .B(new_n188), .C1(KEYINPUT15), .C2(new_n583), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n548), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n192), .A2(G952), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(G234), .B2(G237), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n188), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT21), .B(G898), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n367), .A2(new_n446), .A3(new_n496), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT89), .B(G101), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G3));
  INV_X1    g411(.A(new_n593), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n496), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n582), .B2(new_n583), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT92), .B(G478), .C1(new_n581), .C2(new_n188), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n581), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n578), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n578), .A2(new_n605), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(KEYINPUT33), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n583), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n601), .A2(new_n602), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n543), .B1(new_n542), .B2(new_n532), .ZN(new_n613));
  AOI211_X1 g427(.A(KEYINPUT20), .B(new_n533), .C1(new_n540), .C2(new_n541), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n539), .A2(new_n520), .ZN(new_n615));
  INV_X1    g429(.A(new_n498), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n617), .B2(new_n540), .ZN(new_n618));
  INV_X1    g432(.A(G475), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n613), .A2(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n599), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n330), .A2(new_n340), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n342), .A2(KEYINPUT90), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n188), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n624), .B1(new_n344), .B2(G902), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n626), .A2(new_n627), .A3(new_n242), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n444), .B1(new_n436), .B2(new_n441), .ZN(new_n629));
  AOI211_X1 g443(.A(KEYINPUT79), .B(new_n440), .C1(new_n432), .C2(new_n435), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n622), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n585), .A2(new_n586), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n548), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n599), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n628), .B(new_n636), .C1(new_n629), .C2(new_n630), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  OAI21_X1  g454(.A(KEYINPUT94), .B1(new_n225), .B2(new_n228), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n231), .A2(new_n642), .A3(new_n232), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n641), .B2(new_n643), .ZN(new_n646));
  INV_X1    g460(.A(new_n240), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n238), .A2(new_n648), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n620), .A2(new_n649), .A3(new_n634), .A4(new_n593), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n650), .A2(new_n626), .A3(new_n627), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n496), .C1(new_n629), .C2(new_n630), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(new_n496), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n649), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n629), .B2(new_n630), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n623), .A2(new_n342), .A3(new_n188), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n345), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n341), .A2(KEYINPUT32), .A3(new_n342), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n366), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n591), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n590), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n635), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT95), .B(G128), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G30));
  XNOR2_X1  g485(.A(new_n665), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n446), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT97), .Z(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n676));
  OR3_X1    g490(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT98), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT98), .B1(new_n675), .B2(new_n676), .ZN(new_n678));
  INV_X1    g492(.A(new_n326), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n321), .B1(new_n359), .B2(new_n311), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n188), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n347), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n493), .A2(new_n495), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n620), .A2(new_n447), .A3(new_n649), .A4(new_n634), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n677), .A2(new_n678), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n280), .ZN(G45));
  NOR2_X1   g505(.A1(new_n621), .A2(new_n666), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n661), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n657), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n209), .ZN(G48));
  INV_X1    g509(.A(new_n419), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n412), .B2(new_n414), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n423), .B(KEYINPUT12), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n412), .A2(new_n696), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n698), .B1(new_n699), .B2(KEYINPUT78), .ZN(new_n700));
  INV_X1    g514(.A(new_n429), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n702), .B2(G902), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n441), .A3(new_n432), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(KEYINPUT99), .A3(new_n441), .A4(new_n432), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n367), .A2(new_n622), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND4_X1  g524(.A1(new_n367), .A2(new_n636), .A3(new_n706), .A4(new_n707), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AND2_X1   g526(.A1(new_n703), .A2(new_n432), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n441), .A3(new_n496), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n661), .A3(new_n650), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  OAI21_X1  g531(.A(G472), .B1(new_n344), .B2(G902), .ZN(new_n718));
  NOR2_X1   g532(.A1(G472), .A2(G902), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n328), .A2(new_n329), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n362), .A2(new_n321), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(new_n722), .A3(new_n242), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT100), .B1(new_n548), .B2(new_n587), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n620), .A2(new_n725), .A3(new_n634), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(new_n496), .A3(new_n598), .A4(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n706), .A3(new_n707), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n728), .A2(new_n706), .A3(KEYINPUT101), .A4(new_n707), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n550), .ZN(G24));
  AND2_X1   g548(.A1(new_n718), .A2(new_n722), .ZN(new_n735));
  INV_X1    g549(.A(new_n649), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n692), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n714), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n213), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n440), .B1(new_n436), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n432), .A2(KEYINPUT102), .A3(new_n435), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n741), .A2(KEYINPUT103), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT103), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n493), .A2(new_n447), .A3(new_n495), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n367), .A4(new_n692), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n436), .A2(new_n740), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n441), .A3(new_n742), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT103), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n741), .A2(KEYINPUT103), .A3(new_n742), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n367), .A3(new_n692), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n667), .B(KEYINPUT104), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n746), .A2(new_n758), .A3(new_n367), .A4(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n751), .A2(new_n367), .A3(new_n752), .A4(new_n759), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  OR2_X1    g578(.A1(new_n434), .A2(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n434), .A2(KEYINPUT45), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(G469), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(G469), .A2(G902), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n432), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n768), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n440), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n672), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n612), .A2(new_n548), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT43), .B1(new_n548), .B2(KEYINPUT106), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n775), .B(new_n776), .Z(new_n777));
  AOI21_X1  g591(.A(new_n649), .B1(new_n626), .B2(new_n627), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT44), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT44), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n745), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  XNOR2_X1  g597(.A(new_n773), .B(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n745), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n692), .A2(new_n243), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n661), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  AOI21_X1  g603(.A(new_n784), .B1(new_n440), .B2(new_n713), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n777), .A2(new_n590), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n242), .A3(new_n735), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n790), .A2(new_n745), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n687), .A2(new_n448), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n792), .A2(new_n704), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n735), .A2(new_n736), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n704), .A2(new_n745), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n795), .A2(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n795), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n684), .A2(new_n242), .A3(new_n590), .A4(new_n799), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT114), .Z(new_n806));
  NOR2_X1   g620(.A1(new_n612), .A2(new_n620), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n793), .B(new_n804), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n792), .A2(new_n714), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n813));
  NOR2_X1   g627(.A1(KEYINPUT115), .A2(G953), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n589), .B2(KEYINPUT115), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n801), .A2(new_n367), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT48), .Z(new_n818));
  INV_X1    g632(.A(new_n621), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n816), .B(new_n818), .C1(new_n819), .C2(new_n806), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n637), .A2(new_n652), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n595), .A3(new_n823), .A4(new_n631), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n661), .A2(new_n242), .A3(new_n594), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n496), .B1(new_n629), .B2(new_n630), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n631), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n637), .A2(new_n652), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT107), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n708), .A2(new_n711), .A3(new_n716), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n733), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n749), .A2(new_n750), .ZN(new_n833));
  INV_X1    g647(.A(new_n737), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n752), .A4(new_n785), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n745), .A2(new_n588), .A3(new_n649), .A4(new_n666), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n446), .A2(new_n661), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n830), .A2(new_n832), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n756), .A2(new_n763), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n669), .A2(new_n738), .ZN(new_n843));
  INV_X1    g657(.A(new_n694), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n736), .A2(new_n666), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n741), .A2(new_n742), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n724), .A2(new_n496), .A3(new_n726), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n741), .A2(KEYINPUT108), .A3(new_n742), .A4(new_n845), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n848), .A2(new_n683), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n844), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n669), .A2(new_n694), .A3(new_n738), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n851), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT109), .B1(new_n852), .B2(KEYINPUT110), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n853), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n853), .B1(new_n852), .B2(KEYINPUT109), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT110), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n855), .B2(new_n851), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(KEYINPUT109), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n842), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n858), .B1(new_n865), .B2(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n831), .A2(new_n733), .A3(new_n838), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n756), .A3(new_n763), .A4(new_n830), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(new_n855), .B2(new_n851), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT52), .A2(new_n843), .A3(new_n844), .A4(new_n851), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n868), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT111), .ZN(new_n875));
  XOR2_X1   g689(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n876));
  NAND4_X1  g690(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n860), .A4(new_n864), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n878), .B(new_n868), .C1(new_n870), .C2(new_n873), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n821), .A2(new_n881), .B1(G952), .B2(G953), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n441), .A2(new_n775), .A3(new_n447), .A4(new_n242), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n684), .A2(new_n687), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n713), .B(KEYINPUT49), .Z(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n192), .A2(G952), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(new_n877), .A3(new_n879), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G902), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(G210), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n469), .A2(new_n476), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n474), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT55), .Z(new_n896));
  AOI21_X1  g710(.A(new_n887), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n890), .A2(KEYINPUT117), .A3(G210), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n897), .A2(new_n902), .ZN(G51));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n889), .A2(new_n767), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n876), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n877), .A2(new_n879), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n756), .A2(new_n763), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n857), .A3(new_n830), .A4(new_n869), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n878), .B1(new_n910), .B2(new_n868), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n880), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n768), .B(KEYINPUT57), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n702), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n914), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n912), .B2(new_n880), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT118), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n906), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n904), .B1(new_n921), .B2(new_n887), .ZN(new_n922));
  INV_X1    g736(.A(new_n920), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n430), .B1(new_n919), .B2(KEYINPUT118), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n905), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n887), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n531), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n531), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n887), .ZN(G60));
  INV_X1    g746(.A(new_n609), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n881), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n913), .A2(new_n933), .A3(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n887), .ZN(G63));
  NOR2_X1   g752(.A1(new_n645), .A2(new_n646), .ZN(new_n939));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n888), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT120), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n888), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n229), .A2(new_n233), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n887), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n592), .B2(new_n472), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n830), .A2(new_n832), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n894), .B1(G898), .B2(new_n192), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT122), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n952), .B(new_n954), .ZN(G69));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n855), .B(KEYINPUT124), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n690), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n788), .A2(new_n782), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n745), .B1(new_n621), .B2(new_n635), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n674), .A2(new_n367), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n690), .A2(new_n957), .A3(new_n958), .ZN(new_n965));
  AOI21_X1  g779(.A(G953), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n349), .A2(new_n305), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n502), .B(KEYINPUT123), .Z(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n956), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  INV_X1    g785(.A(new_n965), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n972), .A2(new_n959), .A3(new_n963), .ZN(new_n973));
  OAI211_X1 g787(.A(KEYINPUT125), .B(new_n971), .C1(new_n973), .C2(G953), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n774), .A2(new_n367), .A3(new_n849), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n960), .A2(new_n909), .A3(new_n958), .A4(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n192), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n978), .B(new_n969), .C1(new_n662), .C2(new_n192), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n970), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n981), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n970), .A2(new_n974), .A3(new_n983), .A4(new_n979), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n353), .A2(new_n357), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n326), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n887), .B1(new_n866), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n973), .B2(new_n951), .ZN(new_n992));
  INV_X1    g806(.A(new_n352), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n321), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n988), .B1(new_n977), .B2(new_n951), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT127), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n993), .A2(new_n321), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(G57));
endmodule


