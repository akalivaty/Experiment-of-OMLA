//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202));
  NAND2_X1  g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT74), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n209), .A3(new_n204), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n211), .B2(KEYINPUT82), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n210), .A3(new_n208), .ZN(new_n214));
  INV_X1    g013(.A(new_n207), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT82), .A3(new_n211), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT3), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(G155gat), .B2(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT77), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G155gat), .B(G162gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n221), .A3(new_n222), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(KEYINPUT77), .A3(new_n227), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT29), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n211), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n218), .A2(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n237), .B2(new_n202), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n232), .A2(KEYINPUT77), .A3(new_n227), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n227), .B1(new_n232), .B2(KEYINPUT77), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n235), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n202), .ZN(new_n245));
  INV_X1    g044(.A(new_n237), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n239), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n238), .A2(new_n239), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT83), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G50gat), .ZN(new_n252));
  XOR2_X1   g051(.A(G78gat), .B(G106gat), .Z(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n249), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n248), .A2(new_n249), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n248), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G22gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n256), .A3(new_n262), .A4(new_n254), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G226gat), .ZN(new_n265));
  INV_X1    g064(.A(G233gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT29), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n271), .A2(new_n272), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT23), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(KEYINPUT65), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G169gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT65), .B(G169gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .A3(new_n280), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n278), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n272), .B(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n271), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n275), .B2(new_n279), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n304), .B2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n300), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n303), .A2(new_n305), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n275), .A2(new_n314), .A3(new_n276), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n270), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n268), .B1(new_n299), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n289), .A2(new_n290), .B1(new_n293), .B2(new_n297), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n317), .B1(new_n310), .B2(new_n312), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n321), .A2(new_n267), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n246), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n267), .ZN(new_n325));
  INV_X1    g124(.A(new_n290), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT66), .B1(new_n287), .B2(new_n280), .ZN(new_n327));
  AND4_X1   g126(.A1(KEYINPUT66), .A2(new_n280), .A3(new_n281), .A4(new_n283), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(new_n278), .ZN(new_n330));
  INV_X1    g129(.A(new_n298), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n325), .B(new_n319), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n268), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n321), .B2(new_n322), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n334), .A3(new_n237), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n324), .A2(KEYINPUT75), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n237), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT30), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(KEYINPUT76), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n347), .B1(new_n336), .B2(new_n339), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT30), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n229), .A2(KEYINPUT3), .A3(new_n233), .ZN(new_n353));
  XOR2_X1   g152(.A(G127gat), .B(G134gat), .Z(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(G113gat), .B2(G120gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n354), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT69), .B(G120gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n355), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n244), .A2(new_n353), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n360), .B(new_n364), .C1(new_n242), .C2(new_n243), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n360), .A2(new_n364), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT4), .B1(new_n234), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT79), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n376));
  INV_X1    g175(.A(new_n371), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n234), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n370), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n376), .B(new_n378), .C1(new_n379), .C2(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n369), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n371), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n234), .A2(new_n373), .A3(KEYINPUT4), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n366), .A2(new_n382), .A3(new_n368), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n229), .A3(new_n233), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n368), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n367), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n381), .B2(new_n389), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n389), .A3(new_n394), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n398), .A2(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n264), .B1(new_n352), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n263), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n261), .A2(new_n256), .B1(new_n250), .B2(new_n254), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n395), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n402), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n399), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT80), .B1(new_n399), .B2(KEYINPUT6), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n411), .B(new_n344), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n324), .A2(new_n335), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT38), .B1(new_n415), .B2(KEYINPUT37), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT75), .B(new_n237), .C1(new_n332), .C2(new_n334), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n332), .A2(new_n334), .A3(new_n237), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n337), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n419), .B2(KEYINPUT75), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n347), .B(new_n416), .C1(new_n420), .C2(KEYINPUT37), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT38), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(KEYINPUT37), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n347), .A2(KEYINPUT37), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n348), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n408), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n346), .A2(new_n348), .A3(new_n351), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n375), .A2(new_n380), .A3(new_n366), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n387), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n394), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n370), .A2(new_n385), .A3(new_n368), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT39), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n433), .B2(new_n387), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n432), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(KEYINPUT40), .A3(new_n394), .A4(new_n435), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n431), .A2(new_n409), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n405), .B1(new_n430), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n299), .A2(new_n373), .A3(new_n319), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT70), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n322), .B1(new_n291), .B2(new_n298), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n373), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT71), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n447), .B2(new_n373), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT71), .B(new_n365), .C1(new_n321), .C2(new_n322), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT34), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n450), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT72), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n454), .ZN(new_n459));
  INV_X1    g258(.A(new_n456), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT34), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n446), .A2(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT72), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n455), .A4(new_n456), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT32), .B1(new_n462), .B2(new_n456), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n462), .B2(new_n456), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  OAI221_X1 g272(.A(KEYINPUT32), .B1(new_n467), .B2(new_n473), .C1(new_n462), .C2(new_n456), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n465), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n458), .A2(new_n461), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n474), .A4(new_n464), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT73), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(new_n465), .C1(new_n472), .C2(new_n475), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT36), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n480), .A2(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n406), .B2(new_n407), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n489), .A2(new_n431), .A3(new_n403), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n352), .A2(new_n404), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n479), .A3(new_n264), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT35), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n444), .A2(new_n486), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  AOI21_X1  g298(.A(G1gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n496), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n249), .A2(G15gat), .ZN(new_n502));
  INV_X1    g301(.A(G15gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G22gat), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n502), .A2(new_n504), .A3(new_n497), .ZN(new_n505));
  INV_X1    g304(.A(G1gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT16), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(G8gat), .B1(new_n500), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n498), .A2(new_n507), .A3(new_n499), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n506), .B1(new_n501), .B2(new_n505), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n520), .A2(KEYINPUT15), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n521), .A2(KEYINPUT15), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n520), .A4(new_n522), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n520), .A2(new_n522), .B1(KEYINPUT15), .B2(new_n521), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT17), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n524), .A2(new_n527), .B1(new_n535), .B2(new_n529), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n510), .B(new_n514), .C1(new_n539), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n511), .A2(new_n513), .A3(new_n512), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n510), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n537), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n543), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n550), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n546), .A2(new_n547), .A3(new_n545), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT88), .B1(new_n510), .B2(new_n514), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n540), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n550), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n544), .B(KEYINPUT13), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G197gat), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT11), .B(G169gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n553), .A2(new_n566), .A3(new_n554), .A4(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G64gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G57gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT90), .B(G57gat), .Z(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n572), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT91), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  INV_X1    g379(.A(G78gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n575), .A2(new_n578), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n586), .A2(KEYINPUT89), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n582), .B1(new_n586), .B2(KEYINPUT89), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n577), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G127gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n555), .A2(new_n556), .B1(new_n591), .B2(new_n590), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  INV_X1    g414(.A(G85gat), .ZN(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n611), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n614), .A2(new_n618), .A3(new_n621), .A4(new_n619), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n610), .B1(new_n629), .B2(new_n540), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT17), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n541), .B1(new_n540), .B2(KEYINPUT86), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n630), .B1(new_n633), .B2(new_n629), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT95), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT92), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(new_n630), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n609), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n629), .B1(new_n539), .B2(new_n542), .ZN(new_n643));
  INV_X1    g442(.A(new_n630), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n636), .ZN(new_n645));
  AND4_X1   g444(.A1(new_n642), .A2(new_n645), .A3(new_n640), .A4(new_n609), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n608), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n640), .A3(new_n642), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT96), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n637), .A2(new_n609), .A3(new_n640), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(new_n607), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n623), .A2(new_n625), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n590), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n626), .A2(new_n627), .B1(new_n585), .B2(new_n589), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n589), .A4(new_n585), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n656), .A2(new_n657), .A3(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(G176gat), .B(G204gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n603), .A2(new_n653), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n495), .A2(new_n571), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n403), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT97), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT98), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n673), .A2(new_n431), .ZN(new_n682));
  AOI211_X1 g481(.A(new_n681), .B(new_n682), .C1(new_n679), .C2(new_n678), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n678), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n682), .B2(G8gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(G1325gat));
  NAND3_X1  g485(.A1(new_n673), .A2(new_n503), .A3(new_n487), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n486), .A2(KEYINPUT100), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n484), .A2(new_n689), .A3(new_n485), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n673), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n687), .B1(new_n692), .B2(new_n503), .ZN(G1326gat));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n408), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT101), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n444), .A2(new_n486), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n491), .A2(new_n494), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n653), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n671), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n603), .A2(new_n571), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n403), .A2(new_n517), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n495), .B2(new_n653), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n408), .B1(new_n431), .B2(new_n403), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n398), .A2(new_n400), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(new_n421), .A3(new_n411), .A4(new_n344), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n264), .B1(new_n713), .B2(new_n428), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n440), .A2(new_n442), .A3(new_n409), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n351), .A2(new_n348), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n346), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n485), .B2(new_n484), .ZN(new_n719));
  INV_X1    g518(.A(new_n493), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n431), .A2(new_n403), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(KEYINPUT35), .B1(new_n487), .B2(new_n490), .ZN(new_n723));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n652), .C1(new_n719), .C2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n710), .A2(new_n724), .A3(new_n403), .A4(new_n702), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G29gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n705), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n708), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1328gat));
  NAND4_X1  g529(.A1(new_n700), .A2(new_n515), .A3(new_n431), .A4(new_n702), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT103), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(KEYINPUT103), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n710), .A2(new_n724), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n431), .A3(new_n702), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G36gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n732), .A2(new_n734), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(KEYINPUT46), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT104), .B(new_n733), .C1(new_n732), .C2(new_n734), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n735), .B(new_n738), .C1(new_n741), .C2(new_n742), .ZN(G1329gat));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  INV_X1    g543(.A(new_n486), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n710), .A2(new_n724), .A3(new_n745), .A4(new_n702), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n487), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(G43gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n700), .A2(new_n702), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n744), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n744), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n710), .A2(new_n724), .A3(new_n691), .A4(new_n702), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(G43gat), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT105), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(G43gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n746), .A2(G43gat), .B1(new_n703), .B2(new_n749), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n758), .B(new_n759), .C1(new_n744), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n755), .A2(new_n761), .ZN(G1330gat));
  NAND4_X1  g561(.A1(new_n710), .A2(new_n724), .A3(new_n408), .A4(new_n702), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n698), .A2(new_n699), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n264), .A2(G50gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n765), .A2(new_n652), .A3(new_n702), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(KEYINPUT48), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n767), .B(KEYINPUT106), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n764), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g572(.A(KEYINPUT107), .B(KEYINPUT48), .C1(new_n770), .C2(new_n764), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(G1331gat));
  NAND4_X1  g574(.A1(new_n603), .A2(new_n571), .A3(new_n653), .A4(new_n701), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n495), .B2(new_n776), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n403), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n574), .ZN(G1332gat));
  XNOR2_X1  g582(.A(new_n352), .B(KEYINPUT109), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n778), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT49), .B(G64gat), .Z(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT110), .ZN(G1333gat));
  NAND3_X1  g588(.A1(new_n778), .A2(new_n780), .A3(new_n487), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT111), .A4(new_n487), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n580), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n781), .A2(G71gat), .A3(new_n691), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n408), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n603), .A2(new_n570), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n671), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n736), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n404), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n804), .B1(new_n700), .B2(KEYINPUT112), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n495), .B2(new_n653), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT51), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT112), .B(new_n652), .C1(new_n719), .C2(new_n723), .ZN(new_n812));
  AND4_X1   g611(.A1(KEYINPUT51), .A2(new_n810), .A3(new_n812), .A4(new_n803), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n701), .A2(new_n616), .A3(new_n403), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n736), .A2(new_n784), .A3(new_n805), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(new_n817), .B2(G92gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n784), .A2(new_n617), .A3(new_n701), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT113), .Z(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n810), .A2(new_n812), .A3(new_n803), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n710), .A2(new_n724), .A3(new_n431), .A4(new_n805), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(G92gat), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT52), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n821), .A2(new_n829), .ZN(G1337gat));
  INV_X1    g629(.A(new_n691), .ZN(new_n831));
  OAI21_X1  g630(.A(G99gat), .B1(new_n806), .B2(new_n831), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n748), .A2(G99gat), .A3(new_n671), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n814), .B2(new_n833), .ZN(G1338gat));
  OR2_X1    g633(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g634(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n264), .A2(G106gat), .A3(new_n671), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT114), .Z(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n824), .B2(new_n825), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n710), .A2(new_n724), .A3(new_n408), .A4(new_n805), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n835), .B(new_n836), .C1(new_n840), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n838), .B1(new_n811), .B2(new_n813), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n842), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(G1339gat));
  INV_X1    g646(.A(new_n603), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n668), .B1(new_n662), .B2(KEYINPUT54), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n658), .A2(G230gat), .A3(G233gat), .A4(new_n659), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n662), .A2(new_n853), .A3(KEYINPUT54), .A4(new_n850), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT55), .B(new_n849), .C1(new_n852), .C2(new_n854), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n670), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n559), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n557), .A2(new_n550), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  INV_X1    g661(.A(new_n550), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n510), .A2(new_n514), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n864), .B1(new_n631), .B2(new_n632), .ZN(new_n865));
  OAI211_X1 g664(.A(G229gat), .B(G233gat), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n557), .A2(new_n867), .A3(new_n550), .A4(new_n860), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n565), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n569), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n569), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n652), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n570), .A2(new_n651), .A3(new_n647), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n859), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n652), .A2(new_n671), .A3(new_n871), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n848), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n672), .A2(new_n570), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n408), .B(new_n748), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n784), .A2(new_n404), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n355), .A3(new_n571), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n404), .B1(new_n879), .B2(new_n880), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n720), .ZN(new_n886));
  INV_X1    g685(.A(new_n784), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n570), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n889), .B2(new_n355), .ZN(G1340gat));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n363), .A3(new_n701), .ZN(new_n891));
  OAI21_X1  g690(.A(G120gat), .B1(new_n883), .B2(new_n671), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1341gat));
  NAND3_X1  g692(.A1(new_n888), .A2(new_n595), .A3(new_n603), .ZN(new_n894));
  OAI21_X1  g693(.A(G127gat), .B1(new_n883), .B2(new_n848), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n653), .A2(new_n431), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n886), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n900));
  OAI21_X1  g699(.A(G134gat), .B1(new_n883), .B2(new_n653), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(KEYINPUT56), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n882), .A2(new_n486), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n879), .A2(new_n880), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n408), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n908), .B(new_n264), .C1(new_n879), .C2(new_n880), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n570), .B(new_n905), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G141gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n691), .A2(new_n264), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n885), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n784), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n219), .A3(new_n570), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT58), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n911), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  NAND3_X1  g719(.A1(new_n914), .A2(new_n220), .A3(new_n701), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n408), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n908), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n906), .A2(KEYINPUT57), .A3(new_n408), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n701), .A3(new_n905), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(G148gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n926), .B2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n921), .B1(new_n928), .B2(new_n929), .ZN(G1345gat));
  NAND2_X1  g729(.A1(new_n925), .A2(new_n905), .ZN(new_n931));
  INV_X1    g730(.A(G155gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n848), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n913), .A2(new_n848), .A3(new_n784), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G155gat), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n931), .B2(new_n653), .ZN(new_n939));
  INV_X1    g738(.A(G162gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n898), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n913), .B2(new_n941), .ZN(G1347gat));
  NAND2_X1  g741(.A1(new_n404), .A2(new_n431), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n881), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n571), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n403), .B1(new_n879), .B2(new_n880), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(new_n720), .A3(new_n784), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n287), .A3(new_n570), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n949), .ZN(G1348gat));
  OAI21_X1  g749(.A(G176gat), .B1(new_n945), .B2(new_n671), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n274), .A3(new_n701), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1349gat));
  OAI21_X1  g752(.A(G183gat), .B1(new_n945), .B2(new_n848), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n948), .A2(new_n311), .A3(new_n603), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g756(.A1(new_n948), .A2(new_n308), .A3(new_n652), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n881), .A2(new_n652), .A3(new_n944), .ZN(new_n959));
  XNOR2_X1  g758(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(G190gat), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n959), .B2(G190gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1351gat));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n688), .A2(new_n408), .A3(new_n690), .A4(new_n784), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n947), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n964), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT124), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n965), .A2(new_n964), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(new_n971), .A3(new_n947), .A4(new_n967), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n570), .A3(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(G197gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n831), .A2(new_n944), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n923), .B2(new_n924), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n571), .A2(new_n974), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n973), .A2(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  XOR2_X1   g777(.A(KEYINPUT125), .B(G204gat), .Z(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n671), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n970), .A2(new_n947), .A3(new_n967), .A4(new_n981), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT62), .Z(new_n983));
  AOI21_X1  g782(.A(KEYINPUT126), .B1(new_n976), .B2(new_n701), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n976), .A2(KEYINPUT126), .A3(new_n701), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n980), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n984), .B2(new_n986), .ZN(G1353gat));
  NOR2_X1   g786(.A1(new_n848), .A2(G211gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n972), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n976), .A2(new_n603), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  NOR2_X1   g792(.A1(new_n653), .A2(G218gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n969), .A2(new_n972), .A3(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(new_n975), .ZN(new_n996));
  OAI211_X1 g795(.A(new_n996), .B(new_n652), .C1(new_n907), .C2(new_n909), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G218gat), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n995), .A2(new_n998), .A3(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1355gat));
endmodule


