

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n751), .A2(n980), .ZN(n752) );
  NOR2_X2 U554 ( .A1(G2105), .A2(n522), .ZN(n886) );
  NOR2_X1 U555 ( .A1(G543), .A2(G651), .ZN(n642) );
  INV_X1 U556 ( .A(KEYINPUT30), .ZN(n681) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NOR2_X1 U558 ( .A1(n631), .A2(G651), .ZN(n634) );
  XOR2_X1 U559 ( .A(KEYINPUT66), .B(n529), .Z(n638) );
  XOR2_X1 U560 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  INV_X1 U561 ( .A(G2105), .ZN(n519) );
  NOR2_X1 U562 ( .A1(G2104), .A2(n519), .ZN(n883) );
  NAND2_X1 U563 ( .A1(n883), .A2(G125), .ZN(n527) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n518), .Z(n887) );
  NAND2_X1 U565 ( .A1(G137), .A2(n887), .ZN(n521) );
  INV_X1 U566 ( .A(G2104), .ZN(n522) );
  NOR2_X1 U567 ( .A1(n522), .A2(n519), .ZN(n882) );
  NAND2_X1 U568 ( .A1(G113), .A2(n882), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n525) );
  NAND2_X1 U570 ( .A1(G101), .A2(n886), .ZN(n523) );
  XNOR2_X1 U571 ( .A(KEYINPUT23), .B(n523), .ZN(n524) );
  NOR2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X2 U574 ( .A(KEYINPUT64), .B(n528), .Z(G160) );
  XNOR2_X1 U575 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U576 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U577 ( .A(G132), .ZN(G219) );
  INV_X1 U578 ( .A(G82), .ZN(G220) );
  INV_X1 U579 ( .A(G57), .ZN(G237) );
  NAND2_X1 U580 ( .A1(G88), .A2(n642), .ZN(n531) );
  INV_X1 U581 ( .A(G651), .ZN(n532) );
  OR2_X1 U582 ( .A1(n532), .A2(n631), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G75), .A2(n638), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n538) );
  NAND2_X1 U585 ( .A1(G50), .A2(n634), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n533), .Z(n635) );
  NAND2_X1 U588 ( .A1(G62), .A2(n635), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U590 ( .A(KEYINPUT81), .B(n536), .Z(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G166) );
  NAND2_X1 U592 ( .A1(G52), .A2(n634), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G64), .A2(n635), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U595 ( .A1(G90), .A2(n642), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G77), .A2(n638), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U599 ( .A1(n545), .A2(n544), .ZN(G171) );
  NAND2_X1 U600 ( .A1(n642), .A2(G89), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G76), .A2(n638), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n549), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U605 ( .A1(G51), .A2(n634), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G63), .A2(n635), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U610 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U613 ( .A(n556), .B(KEYINPUT10), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT68), .B(n557), .ZN(G223) );
  XOR2_X1 U615 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n559) );
  INV_X1 U616 ( .A(G223), .ZN(n821) );
  NAND2_X1 U617 ( .A1(n821), .A2(G567), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT69), .B(n560), .Z(G234) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(KEYINPUT71), .Z(n562) );
  NAND2_X1 U621 ( .A1(G56), .A2(n635), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n562), .B(n561), .ZN(n571) );
  NAND2_X1 U623 ( .A1(G43), .A2(n634), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT72), .B(n563), .Z(n569) );
  NAND2_X1 U625 ( .A1(n642), .A2(G81), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G68), .A2(n638), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X2 U632 ( .A(KEYINPUT73), .B(n572), .ZN(n984) );
  NAND2_X1 U633 ( .A1(G860), .A2(n984), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n573), .B(KEYINPUT74), .ZN(G153) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G92), .A2(n642), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G79), .A2(n638), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G54), .A2(n634), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G66), .A2(n635), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT15), .ZN(n970) );
  INV_X1 U645 ( .A(G868), .ZN(n652) );
  NAND2_X1 U646 ( .A1(n970), .A2(n652), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G53), .A2(n634), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G65), .A2(n635), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G91), .A2(n642), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G78), .A2(n638), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n962) );
  INV_X1 U655 ( .A(n962), .ZN(G299) );
  NOR2_X1 U656 ( .A1(G286), .A2(n652), .ZN(n590) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G297) );
  INV_X1 U659 ( .A(G559), .ZN(n591) );
  NOR2_X1 U660 ( .A1(G860), .A2(n591), .ZN(n592) );
  XNOR2_X1 U661 ( .A(KEYINPUT75), .B(n592), .ZN(n593) );
  INV_X1 U662 ( .A(n970), .ZN(n610) );
  NAND2_X1 U663 ( .A1(n593), .A2(n610), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G559), .A2(n970), .ZN(n595) );
  NOR2_X1 U666 ( .A1(n652), .A2(n595), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n984), .A2(G868), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT76), .B(n598), .Z(G282) );
  XNOR2_X1 U670 ( .A(G2100), .B(KEYINPUT79), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G99), .A2(n886), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G111), .A2(n882), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n887), .A2(G135), .ZN(n601) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(n601), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n883), .A2(G123), .ZN(n602) );
  XOR2_X1 U677 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U679 ( .A(KEYINPUT78), .B(n605), .Z(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n914) );
  XNOR2_X1 U681 ( .A(n914), .B(G2096), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G156) );
  XOR2_X1 U683 ( .A(n984), .B(KEYINPUT80), .Z(n612) );
  NAND2_X1 U684 ( .A1(G559), .A2(n610), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n612), .B(n611), .ZN(n650) );
  NOR2_X1 U686 ( .A1(G860), .A2(n650), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G55), .A2(n634), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G67), .A2(n635), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G93), .A2(n642), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G80), .A2(n638), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n653) );
  XOR2_X1 U694 ( .A(n619), .B(n653), .Z(G145) );
  NAND2_X1 U695 ( .A1(n635), .A2(G60), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G47), .A2(n634), .ZN(n620) );
  XOR2_X1 U697 ( .A(KEYINPUT67), .B(n620), .Z(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G85), .A2(n642), .ZN(n623) );
  XNOR2_X1 U700 ( .A(KEYINPUT65), .B(n623), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G72), .A2(n638), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U704 ( .A1(G49), .A2(n634), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n635), .A2(n630), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G48), .A2(n634), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G61), .A2(n635), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n638), .A2(G73), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U716 ( .A1(n642), .A2(G86), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(G305) );
  XNOR2_X1 U718 ( .A(KEYINPUT19), .B(G290), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(G288), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(n653), .ZN(n648) );
  XNOR2_X1 U721 ( .A(G166), .B(n962), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(G305), .ZN(n849) );
  XOR2_X1 U724 ( .A(n849), .B(n650), .Z(n651) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G868), .A2(n653), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G2072), .A2(n660), .ZN(G158) );
  NAND2_X1 U734 ( .A1(G69), .A2(G120), .ZN(n661) );
  NOR2_X1 U735 ( .A1(G237), .A2(n661), .ZN(n662) );
  NAND2_X1 U736 ( .A1(G108), .A2(n662), .ZN(n904) );
  NAND2_X1 U737 ( .A1(G567), .A2(n904), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT83), .ZN(n668) );
  NOR2_X1 U739 ( .A1(G220), .A2(G219), .ZN(n664) );
  XNOR2_X1 U740 ( .A(KEYINPUT22), .B(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G96), .ZN(n666) );
  OR2_X1 U742 ( .A1(G218), .A2(n666), .ZN(n905) );
  AND2_X1 U743 ( .A1(G2106), .A2(n905), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n668), .A2(n667), .ZN(G319) );
  INV_X1 U745 ( .A(G319), .ZN(n670) );
  NAND2_X1 U746 ( .A1(G483), .A2(G661), .ZN(n669) );
  NOR2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n824) );
  NAND2_X1 U748 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U749 ( .A1(G102), .A2(n886), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G138), .A2(n887), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U752 ( .A1(G114), .A2(n882), .ZN(n674) );
  NAND2_X1 U753 ( .A1(G126), .A2(n883), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n676), .A2(n675), .ZN(G164) );
  INV_X1 U756 ( .A(G166), .ZN(G303) );
  NAND2_X1 U757 ( .A1(G40), .A2(G160), .ZN(n762) );
  INV_X1 U758 ( .A(n762), .ZN(n677) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n763) );
  NAND2_X2 U760 ( .A1(n677), .A2(n763), .ZN(n721) );
  NAND2_X2 U761 ( .A1(G8), .A2(n721), .ZN(n758) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n678) );
  XOR2_X1 U763 ( .A(n678), .B(KEYINPUT24), .Z(n679) );
  NOR2_X1 U764 ( .A1(n758), .A2(n679), .ZN(n753) );
  NOR2_X1 U765 ( .A1(G1966), .A2(n758), .ZN(n733) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n721), .ZN(n730) );
  NOR2_X1 U767 ( .A1(n733), .A2(n730), .ZN(n680) );
  AND2_X1 U768 ( .A1(n680), .A2(G8), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U770 ( .A1(G168), .A2(n683), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n684), .B(KEYINPUT91), .ZN(n688) );
  XOR2_X1 U772 ( .A(G2078), .B(KEYINPUT25), .Z(n941) );
  NOR2_X1 U773 ( .A1(n941), .A2(n721), .ZN(n686) );
  INV_X1 U774 ( .A(n721), .ZN(n696) );
  NOR2_X1 U775 ( .A1(n696), .A2(G1961), .ZN(n685) );
  NOR2_X1 U776 ( .A1(n686), .A2(n685), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n714), .A2(G301), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT31), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n696), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  AND2_X1 U782 ( .A1(G1956), .A2(n721), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n962), .A2(n695), .ZN(n694) );
  XNOR2_X1 U785 ( .A(KEYINPUT89), .B(KEYINPUT28), .ZN(n693) );
  XNOR2_X1 U786 ( .A(n694), .B(n693), .ZN(n712) );
  NAND2_X1 U787 ( .A1(n962), .A2(n695), .ZN(n710) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n721), .ZN(n698) );
  NAND2_X1 U789 ( .A1(G2067), .A2(n696), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n970), .A2(n706), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n984), .A2(n699), .ZN(n705) );
  INV_X1 U793 ( .A(G1996), .ZN(n937) );
  NOR2_X1 U794 ( .A1(n721), .A2(n937), .ZN(n701) );
  XOR2_X1 U795 ( .A(KEYINPUT26), .B(KEYINPUT90), .Z(n700) );
  XNOR2_X1 U796 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n721), .A2(G1341), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n706), .A2(n970), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U804 ( .A(KEYINPUT29), .B(n713), .Z(n717) );
  NOR2_X1 U805 ( .A1(n714), .A2(G301), .ZN(n715) );
  XOR2_X1 U806 ( .A(KEYINPUT88), .B(n715), .Z(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U809 ( .A(n720), .B(KEYINPUT92), .ZN(n731) );
  NAND2_X1 U810 ( .A1(n731), .A2(G286), .ZN(n728) );
  INV_X1 U811 ( .A(G8), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n758), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n721), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U818 ( .A(n729), .B(KEYINPUT32), .ZN(n737) );
  NAND2_X1 U819 ( .A1(G8), .A2(n730), .ZN(n735) );
  INV_X1 U820 ( .A(n731), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n756) );
  INV_X1 U824 ( .A(G1971), .ZN(n1005) );
  NAND2_X1 U825 ( .A1(G166), .A2(n1005), .ZN(n960) );
  INV_X1 U826 ( .A(n960), .ZN(n738) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NOR2_X1 U828 ( .A1(n738), .A2(n965), .ZN(n739) );
  AND2_X1 U829 ( .A1(n756), .A2(n739), .ZN(n740) );
  NOR2_X1 U830 ( .A1(n758), .A2(n740), .ZN(n745) );
  NAND2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n968) );
  INV_X1 U832 ( .A(KEYINPUT33), .ZN(n747) );
  INV_X1 U833 ( .A(n758), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n741), .A2(n965), .ZN(n742) );
  NOR2_X1 U835 ( .A1(n747), .A2(n742), .ZN(n743) );
  XNOR2_X1 U836 ( .A(n743), .B(KEYINPUT93), .ZN(n746) );
  AND2_X1 U837 ( .A1(n968), .A2(n746), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n750) );
  INV_X1 U839 ( .A(n746), .ZN(n748) );
  OR2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n749) );
  AND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U842 ( .A(G1981), .B(G305), .ZN(n980) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n761) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U845 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT94), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n794) );
  NOR2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n806) );
  XNOR2_X1 U851 ( .A(G2067), .B(KEYINPUT37), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(KEYINPUT84), .ZN(n804) );
  NAND2_X1 U853 ( .A1(G104), .A2(n886), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G140), .A2(n887), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U856 ( .A(KEYINPUT34), .B(n767), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G116), .A2(n882), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G128), .A2(n883), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U860 ( .A(KEYINPUT35), .B(n770), .Z(n771) );
  NOR2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT36), .B(n773), .ZN(n871) );
  NOR2_X1 U863 ( .A1(n804), .A2(n871), .ZN(n918) );
  NAND2_X1 U864 ( .A1(n806), .A2(n918), .ZN(n801) );
  XNOR2_X1 U865 ( .A(G1986), .B(G290), .ZN(n959) );
  AND2_X1 U866 ( .A1(n959), .A2(n806), .ZN(n791) );
  XNOR2_X1 U867 ( .A(n806), .B(KEYINPUT86), .ZN(n789) );
  NAND2_X1 U868 ( .A1(G141), .A2(n887), .ZN(n775) );
  NAND2_X1 U869 ( .A1(G117), .A2(n882), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n886), .A2(G105), .ZN(n776) );
  XOR2_X1 U872 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n883), .A2(G129), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n861) );
  NAND2_X1 U876 ( .A1(G1996), .A2(n861), .ZN(n788) );
  XOR2_X1 U877 ( .A(KEYINPUT85), .B(G1991), .Z(n934) );
  NAND2_X1 U878 ( .A1(G95), .A2(n886), .ZN(n782) );
  NAND2_X1 U879 ( .A1(G107), .A2(n882), .ZN(n781) );
  NAND2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U881 ( .A1(G131), .A2(n887), .ZN(n784) );
  NAND2_X1 U882 ( .A1(G119), .A2(n883), .ZN(n783) );
  NAND2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n869) );
  NAND2_X1 U885 ( .A1(n934), .A2(n869), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n788), .A2(n787), .ZN(n912) );
  NAND2_X1 U887 ( .A1(n789), .A2(n912), .ZN(n790) );
  XNOR2_X1 U888 ( .A(n790), .B(KEYINPUT87), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n791), .A2(n798), .ZN(n792) );
  AND2_X1 U890 ( .A1(n801), .A2(n792), .ZN(n793) );
  NAND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n809) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n861), .ZN(n908) );
  NOR2_X1 U893 ( .A1(n934), .A2(n869), .ZN(n915) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n795) );
  NOR2_X1 U895 ( .A1(n915), .A2(n795), .ZN(n796) );
  XOR2_X1 U896 ( .A(KEYINPUT95), .B(n796), .Z(n797) );
  NOR2_X1 U897 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U898 ( .A1(n908), .A2(n799), .ZN(n800) );
  XNOR2_X1 U899 ( .A(n800), .B(KEYINPUT39), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U901 ( .A(n803), .B(KEYINPUT96), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n804), .A2(n871), .ZN(n911) );
  NAND2_X1 U903 ( .A1(n805), .A2(n911), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n810), .ZN(G329) );
  XOR2_X1 U907 ( .A(KEYINPUT97), .B(G2427), .Z(n812) );
  XNOR2_X1 U908 ( .A(G2435), .B(G2438), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n812), .B(n811), .ZN(n819) );
  XOR2_X1 U910 ( .A(G2443), .B(G2430), .Z(n814) );
  XNOR2_X1 U911 ( .A(G2454), .B(G2446), .ZN(n813) );
  XNOR2_X1 U912 ( .A(n814), .B(n813), .ZN(n815) );
  XOR2_X1 U913 ( .A(n815), .B(G2451), .Z(n817) );
  XNOR2_X1 U914 ( .A(G1348), .B(G1341), .ZN(n816) );
  XNOR2_X1 U915 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n820), .A2(G14), .ZN(n898) );
  XOR2_X1 U918 ( .A(KEYINPUT98), .B(n898), .Z(G401) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U921 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U923 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n826) );
  XNOR2_X1 U925 ( .A(KEYINPUT42), .B(G2678), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U927 ( .A(KEYINPUT100), .B(G2090), .Z(n828) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U931 ( .A(G2100), .B(G2096), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n834) );
  XOR2_X1 U933 ( .A(G2078), .B(G2084), .Z(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1971), .B(G1976), .Z(n836) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n846) );
  XOR2_X1 U938 ( .A(KEYINPUT102), .B(KEYINPUT41), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1981), .B(KEYINPUT103), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U941 ( .A(G1961), .B(G1956), .Z(n840) );
  XNOR2_X1 U942 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U945 ( .A(KEYINPUT104), .B(G2474), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(G229) );
  XNOR2_X1 U948 ( .A(G286), .B(KEYINPUT111), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n970), .B(G171), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n851) );
  XOR2_X1 U951 ( .A(n984), .B(n849), .Z(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  NOR2_X1 U953 ( .A1(G37), .A2(n852), .ZN(G397) );
  NAND2_X1 U954 ( .A1(G124), .A2(n883), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G136), .A2(n887), .ZN(n854) );
  XOR2_X1 U957 ( .A(KEYINPUT105), .B(n854), .Z(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G100), .A2(n886), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G112), .A2(n882), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  XNOR2_X1 U963 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n861), .B(KEYINPUT46), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(KEYINPUT106), .B(n864), .ZN(n866) );
  XNOR2_X1 U967 ( .A(G160), .B(KEYINPUT48), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U969 ( .A(G164), .B(n867), .Z(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n914), .B(n870), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n871), .B(G162), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n895) );
  NAND2_X1 U974 ( .A1(G103), .A2(n886), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G139), .A2(n887), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n883), .A2(G127), .ZN(n876) );
  XOR2_X1 U978 ( .A(KEYINPUT107), .B(n876), .Z(n878) );
  NAND2_X1 U979 ( .A1(n882), .A2(G115), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n923) );
  NAND2_X1 U983 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n923), .B(n893), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U994 ( .A(KEYINPUT110), .B(n897), .ZN(G395) );
  NAND2_X1 U995 ( .A1(G319), .A2(n898), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(n899), .ZN(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G397), .A2(G395), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(G225) );
  XOR2_X1 U1001 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  INV_X1 U1003 ( .A(G120), .ZN(G236) );
  INV_X1 U1004 ( .A(G96), .ZN(G221) );
  INV_X1 U1005 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(KEYINPUT99), .B(n906), .ZN(G261) );
  INV_X1 U1008 ( .A(G261), .ZN(G325) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1010 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1012 ( .A(KEYINPUT114), .B(n909), .Z(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT51), .B(n910), .ZN(n931) );
  INV_X1 U1014 ( .A(n911), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(G2084), .B(G160), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT113), .B(n920), .Z(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G2072), .B(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n926), .Z(n927) );
  XNOR2_X1 U1026 ( .A(KEYINPUT115), .B(n927), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n932), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1031 ( .A(n934), .B(G25), .ZN(n946) );
  XNOR2_X1 U1032 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G32), .B(KEYINPUT116), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G27), .B(n941), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(G28), .A2(n947), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n948), .ZN(n952) );
  XOR2_X1 U1044 ( .A(G34), .B(KEYINPUT118), .Z(n950) );
  XNOR2_X1 U1045 ( .A(G2084), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(n950), .B(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(KEYINPUT119), .B(n955), .Z(n956) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n956), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT55), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G11), .ZN(n1020) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .ZN(n989) );
  INV_X1 U1055 ( .A(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n977) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n975) );
  XNOR2_X1 U1058 ( .A(G1956), .B(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1061 ( .A(n965), .B(KEYINPUT121), .Z(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n970), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT120), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT122), .B(n978), .Z(n983) );
  XOR2_X1 U1070 ( .A(G1966), .B(G168), .Z(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT57), .B(n981), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n987) );
  XOR2_X1 U1074 ( .A(n984), .B(G1341), .Z(n985) );
  XNOR2_X1 U1075 ( .A(KEYINPUT123), .B(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n1018) );
  INV_X1 U1078 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1079 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n1000) );
  XNOR2_X1 U1080 ( .A(KEYINPUT59), .B(G1348), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(G4), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(G1956), .B(G20), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT124), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G19), .B(G1341), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n994), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n1000), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G5), .B(G1961), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(G22), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G1986), .B(G24), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G1976), .B(G23), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

