//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n197), .C1(G119), .C2(new_n196), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT24), .B(G110), .Z(new_n200));
  XNOR2_X1  g014(.A(G119), .B(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n192), .A2(new_n203), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n198), .A2(G110), .B1(new_n201), .B2(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n190), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(new_n189), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(G146), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(KEYINPUT22), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(G137), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G902), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n208), .A3(new_n213), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G234), .ZN(new_n221));
  OAI21_X1  g035(.A(G217), .B1(new_n221), .B2(G902), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT74), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(KEYINPUT75), .A3(new_n224), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n218), .A2(new_n224), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n232));
  INV_X1    g046(.A(G134), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(G137), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(G137), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n234), .A2(new_n237), .A3(new_n240), .A4(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT64), .B(G143), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n246), .B(new_n247), .C1(new_n248), .C2(G146), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT64), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT64), .A2(G143), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n191), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n191), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n244), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n250), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT64), .A2(G143), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT64), .A2(G143), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(G146), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n254), .ZN(new_n262));
  OAI21_X1  g076(.A(G146), .B1(new_n259), .B2(new_n260), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n191), .A2(G143), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(KEYINPUT0), .A3(G128), .A4(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n243), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n236), .A2(G134), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n233), .A2(G137), .ZN(new_n269));
  OAI21_X1  g083(.A(G131), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n241), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n263), .A2(new_n264), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n263), .A2(new_n275), .A3(new_n264), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n253), .A2(new_n255), .B1(new_n278), .B2(G128), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n271), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n282));
  INV_X1    g096(.A(G113), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT67), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(KEYINPUT2), .B2(G113), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n284), .A2(new_n286), .B1(KEYINPUT2), .B2(G113), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n194), .A2(KEYINPUT68), .A3(G116), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  INV_X1    g104(.A(G116), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(G119), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT69), .B(G116), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n289), .B(new_n292), .C1(new_n293), .C2(new_n194), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G116), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n287), .A2(new_n300), .A3(new_n289), .A4(new_n292), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n267), .A2(new_n281), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT28), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n249), .A2(new_n256), .A3(new_n244), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT70), .B1(new_n262), .B2(new_n265), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n242), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n246), .B1(new_n248), .B2(G146), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n275), .B1(new_n309), .B2(new_n272), .ZN(new_n310));
  INV_X1    g124(.A(new_n276), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n280), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n271), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n302), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n308), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT71), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(G101), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n210), .A3(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(KEYINPUT29), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n302), .B1(new_n267), .B2(new_n281), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n327), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT72), .B1(new_n327), .B2(KEYINPUT28), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n319), .B(new_n325), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n216), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT73), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n333), .A3(new_n216), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n308), .A2(new_n314), .A3(KEYINPUT30), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n242), .A2(new_n265), .A3(new_n262), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n279), .B1(new_n274), .B2(new_n276), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n271), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n241), .A2(new_n270), .A3(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT30), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n344), .A3(new_n302), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n316), .ZN(new_n346));
  INV_X1    g160(.A(new_n324), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n340), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT65), .B1(new_n241), .B2(new_n270), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n312), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n315), .B1(new_n352), .B2(new_n336), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT28), .B1(new_n303), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n304), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n316), .A2(KEYINPUT71), .A3(new_n317), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n348), .B1(new_n347), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n332), .A2(new_n334), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G472), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n345), .A2(new_n324), .A3(new_n316), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n345), .A2(KEYINPUT31), .A3(new_n324), .A4(new_n316), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n347), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n363), .A2(new_n364), .B1(new_n357), .B2(new_n347), .ZN(new_n371));
  INV_X1    g185(.A(new_n369), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT32), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n231), .B1(new_n360), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n383), .B(KEYINPUT3), .C1(new_n376), .C2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n378), .A2(new_n379), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n382), .A2(new_n379), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n378), .A4(new_n384), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(G101), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n392), .C1(new_n306), .C2(new_n307), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n257), .A2(new_n266), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(KEYINPUT78), .A3(new_n392), .A4(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n309), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n400));
  OAI21_X1  g214(.A(G128), .B1(new_n261), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n277), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  INV_X1    g218(.A(new_n379), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n376), .A2(G107), .ZN(new_n406));
  OAI21_X1  g220(.A(G101), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n389), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n389), .A2(new_n407), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT10), .B1(new_n337), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n398), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n242), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n398), .A2(new_n243), .A3(new_n412), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n210), .A2(G227), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n416), .B(new_n417), .Z(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n418), .ZN(new_n420));
  AOI221_X4 g234(.A(new_n242), .B1(new_n409), .B2(new_n411), .C1(new_n395), .C2(new_n397), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n277), .A2(new_n410), .A3(new_n280), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n274), .A2(new_n276), .B1(new_n399), .B2(new_n401), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n424), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT12), .B1(new_n424), .B2(new_n242), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n420), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(new_n428), .A3(G469), .ZN(new_n429));
  NAND2_X1  g243(.A1(G469), .A2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT79), .B1(new_n421), .B2(new_n420), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n425), .A2(new_n426), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n415), .A2(new_n434), .A3(new_n418), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n243), .B1(new_n398), .B2(new_n412), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n420), .B1(new_n421), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(G902), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n431), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n210), .A2(G952), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G234), .B2(G237), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT21), .B(G898), .Z(new_n445));
  OAI211_X1 g259(.A(G902), .B(G953), .C1(new_n221), .C2(new_n322), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT90), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n187), .B(new_n280), .C1(new_n310), .C2(new_n311), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n210), .A2(G224), .ZN(new_n453));
  OAI21_X1  g267(.A(G125), .B1(new_n249), .B2(new_n256), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(KEYINPUT7), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n389), .A2(new_n458), .A3(new_n407), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT82), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n194), .A3(G116), .ZN(new_n462));
  OAI211_X1 g276(.A(G113), .B(new_n462), .C1(new_n294), .C2(new_n461), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n301), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n460), .B(new_n464), .C1(KEYINPUT82), .C2(new_n410), .ZN(new_n465));
  XOR2_X1   g279(.A(G110), .B(G122), .Z(new_n466));
  XOR2_X1   g280(.A(new_n466), .B(KEYINPUT8), .Z(new_n467));
  NAND4_X1  g281(.A1(new_n459), .A2(new_n463), .A3(KEYINPUT82), .A4(new_n301), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(KEYINPUT83), .A3(new_n467), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n452), .A2(new_n454), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(KEYINPUT7), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n390), .A2(new_n302), .A3(new_n392), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n408), .A2(new_n301), .A3(new_n463), .ZN(new_n477));
  INV_X1    g291(.A(new_n466), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n457), .A2(new_n471), .A3(new_n472), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n466), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n484));
  INV_X1    g298(.A(new_n453), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n473), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n487), .A3(new_n466), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n216), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n492), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n481), .A2(new_n216), .A3(new_n489), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n451), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n296), .B2(new_n298), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n291), .A2(G122), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n504), .B(G107), .C1(new_n501), .C2(new_n500), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n381), .B(new_n503), .C1(new_n293), .C2(new_n498), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n245), .A2(G128), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n248), .B2(G128), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n233), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G107), .B1(new_n499), .B2(new_n502), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n511), .A2(new_n506), .B1(new_n233), .B2(new_n508), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n248), .A2(new_n514), .A3(G128), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n259), .A2(new_n260), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n196), .ZN(new_n518));
  OAI211_X1 g332(.A(G134), .B(new_n515), .C1(new_n518), .C2(new_n514), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n512), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n513), .B1(new_n512), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT9), .B(G234), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(G217), .A3(new_n210), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n510), .B(new_n526), .C1(new_n520), .C2(new_n521), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n527), .ZN(new_n528));
  OR3_X1    g342(.A1(new_n522), .A2(KEYINPUT88), .A3(new_n524), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n216), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n529), .A3(new_n216), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n523), .ZN(new_n540));
  OAI21_X1  g354(.A(G221), .B1(new_n540), .B2(G902), .ZN(new_n541));
  XOR2_X1   g355(.A(new_n541), .B(KEYINPUT76), .Z(new_n542));
  NOR4_X1   g356(.A1(new_n441), .A2(new_n497), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G475), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n322), .A2(new_n210), .A3(G214), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n517), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n245), .A2(new_n322), .A3(new_n210), .A4(G214), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n240), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(G131), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(new_n550), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n192), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G113), .B(G122), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n376), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n546), .A2(KEYINPUT18), .A3(G131), .A4(new_n547), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n189), .B(new_n191), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n558), .A2(new_n549), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n554), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n549), .A2(new_n551), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n207), .A2(KEYINPUT19), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n189), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n191), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n206), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n568), .B2(new_n561), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n544), .B(new_n216), .C1(new_n562), .C2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n569), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n554), .A2(new_n556), .A3(new_n561), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(KEYINPUT20), .A3(new_n544), .A4(new_n216), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT86), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n554), .A2(new_n561), .ZN(new_n579));
  INV_X1    g393(.A(new_n556), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(KEYINPUT86), .B(new_n556), .C1(new_n554), .C2(new_n561), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n544), .B1(new_n583), .B2(new_n216), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n375), .A2(new_n543), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND2_X1  g401(.A1(new_n530), .A2(new_n531), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n528), .A2(new_n529), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n525), .A2(KEYINPUT33), .A3(new_n527), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(G478), .A3(new_n216), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n585), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n449), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n493), .B2(new_n495), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n448), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT91), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n367), .A2(new_n216), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n367), .A2(new_n369), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR4_X1   g415(.A1(new_n601), .A2(new_n441), .A3(new_n231), .A4(new_n542), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G104), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n603), .B(new_n605), .ZN(G6));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n448), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n539), .A2(new_n585), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NAND2_X1  g426(.A1(new_n227), .A2(new_n228), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n214), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n209), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n216), .A3(new_n223), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT93), .Z(new_n617));
  NOR2_X1   g431(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n601), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n543), .A2(new_n585), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT37), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(G110), .Z(G12));
  INV_X1    g436(.A(new_n595), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n360), .B2(new_n374), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n436), .A2(new_n438), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n440), .A3(new_n216), .ZN(new_n626));
  INV_X1    g440(.A(new_n431), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n542), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n618), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n443), .B(KEYINPUT94), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(G900), .B2(new_n446), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT95), .Z(new_n633));
  NOR2_X1   g447(.A1(new_n608), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n624), .A2(new_n628), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G128), .ZN(G30));
  XOR2_X1   g450(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n493), .A2(new_n639), .A3(new_n495), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n639), .B1(new_n493), .B2(new_n495), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n493), .A2(new_n495), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n493), .A2(new_n639), .A3(new_n495), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n539), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n585), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n633), .B(KEYINPUT39), .Z(new_n652));
  AND2_X1   g466(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n655), .A3(new_n449), .A4(new_n618), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  INV_X1    g471(.A(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n327), .A2(new_n347), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n361), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n361), .A2(KEYINPUT98), .A3(new_n659), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(KEYINPUT99), .B(new_n664), .C1(new_n373), .C2(new_n370), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  INV_X1    g480(.A(new_n664), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n374), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n657), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n371), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n374), .A2(new_n666), .A3(new_n667), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(KEYINPUT100), .A3(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n669), .B(new_n675), .C1(new_n654), .C2(new_n653), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n656), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n248), .ZN(G45));
  NAND2_X1  g492(.A1(new_n592), .A2(new_n588), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n577), .A2(new_n584), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n633), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n624), .A2(new_n628), .A3(new_n629), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  INV_X1    g498(.A(new_n597), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n439), .A2(new_n440), .ZN(new_n686));
  AOI211_X1 g500(.A(G469), .B(G902), .C1(new_n436), .C2(new_n438), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n542), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n375), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT41), .B(G113), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND3_X1  g506(.A1(new_n375), .A2(new_n609), .A3(new_n688), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  AND2_X1   g508(.A1(new_n624), .A2(new_n629), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n688), .A2(new_n585), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n695), .A2(new_n648), .A3(new_n448), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AND2_X1   g513(.A1(new_n688), .A2(new_n649), .ZN(new_n700));
  INV_X1    g514(.A(new_n231), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT101), .B(G472), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n319), .B1(new_n328), .B2(new_n329), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n347), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n365), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n598), .A2(new_n702), .B1(new_n705), .B2(new_n369), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n607), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT102), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n625), .A2(new_n216), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  INV_X1    g527(.A(new_n542), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n595), .A3(new_n714), .A4(new_n626), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n682), .A2(new_n706), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n629), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  NAND2_X1  g533(.A1(new_n441), .A2(KEYINPUT103), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n687), .B2(new_n431), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n493), .A2(new_n495), .A3(new_n449), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n542), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n720), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n375), .A3(new_n682), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n375), .A4(new_n682), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT104), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n240), .ZN(G33));
  NAND3_X1  g546(.A1(new_n725), .A2(new_n375), .A3(new_n634), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n419), .A2(new_n428), .A3(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n419), .B2(new_n428), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n735), .B(G469), .C1(new_n738), .C2(G902), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n419), .A2(new_n428), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n419), .A2(new_n428), .A3(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(G469), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n430), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n626), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n714), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n652), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n679), .A2(new_n585), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n629), .A3(new_n601), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n723), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n748), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NAND2_X1  g571(.A1(new_n360), .A2(new_n374), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n746), .A2(new_n760), .A3(new_n714), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n746), .B2(new_n714), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n746), .A2(new_n714), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n746), .A2(new_n760), .A3(new_n714), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n758), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n723), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n231), .A3(new_n682), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NOR2_X1   g585(.A1(new_n686), .A2(new_n687), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT106), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n542), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n767), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n749), .A2(new_n750), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n679), .B2(new_n585), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n630), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n707), .A3(new_n723), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT112), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n763), .A2(new_n767), .A3(KEYINPUT117), .A4(new_n774), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n686), .A2(new_n687), .A3(new_n542), .A4(new_n449), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n647), .A2(KEYINPUT113), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n780), .A2(new_n707), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n642), .A2(new_n646), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n713), .A2(new_n714), .A3(new_n626), .A4(new_n594), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n669), .A2(new_n675), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n772), .A2(new_n701), .A3(new_n724), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n679), .A2(new_n680), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n443), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n786), .A2(new_n791), .A3(new_n787), .A4(new_n794), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n772), .A2(new_n724), .ZN(new_n803));
  INV_X1    g617(.A(new_n780), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n629), .A4(new_n706), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n803), .A2(new_n804), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n758), .A2(new_n701), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n809), .A2(KEYINPUT48), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT48), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n798), .A2(new_n443), .A3(new_n593), .A4(new_n799), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n442), .B1(new_n787), .B2(new_n716), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n813), .A2(KEYINPUT118), .A3(new_n814), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n808), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n801), .A2(new_n802), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n805), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n797), .B2(new_n806), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n775), .A2(new_n782), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n821), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT119), .ZN(new_n835));
  INV_X1    g649(.A(new_n689), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n836), .A2(new_n597), .B1(new_n708), .B2(new_n700), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT108), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n698), .A4(new_n693), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n709), .B1(new_n685), .B2(new_n689), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n624), .A2(new_n648), .A3(new_n448), .A4(new_n629), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n693), .B1(new_n841), .B2(new_n696), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT108), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n608), .A2(KEYINPUT109), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT109), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n539), .A2(new_n585), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n496), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT110), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n593), .A2(new_n496), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(new_n851), .A3(new_n496), .A4(new_n847), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n602), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n854), .A2(new_n586), .A3(new_n620), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n717), .A2(new_n722), .A3(new_n720), .A4(new_n724), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n723), .A2(new_n633), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n758), .A2(new_n648), .A3(new_n628), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n858), .B2(new_n680), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n629), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n730), .A2(new_n855), .A3(new_n860), .A4(new_n733), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n720), .A2(new_n722), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n673), .A2(new_n674), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n623), .A2(new_n650), .A3(new_n633), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n714), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n629), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n635), .A2(new_n683), .A3(new_n718), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n635), .A2(new_n718), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n720), .A2(new_n722), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n674), .B2(new_n673), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n714), .A3(new_n618), .A4(new_n865), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT52), .A4(new_n683), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n844), .A2(new_n861), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n730), .A2(new_n855), .A3(new_n860), .A4(new_n733), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n843), .B2(new_n839), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n867), .B2(new_n868), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT53), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n877), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n882), .B2(new_n874), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n840), .A2(new_n842), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n861), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n821), .A2(new_n831), .A3(new_n895), .A4(new_n833), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n835), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g711(.A1(G952), .A2(G953), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n773), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n231), .B(new_n542), .C1(new_n900), .C2(KEYINPUT49), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(new_n585), .A3(new_n450), .A4(new_n679), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT107), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n900), .A2(KEYINPUT49), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n798), .A3(new_n647), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(G75));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n887), .A2(new_n891), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G902), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n494), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n484), .A2(new_n488), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n486), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n910), .A2(new_n915), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n210), .A2(G952), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G51));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n879), .B2(new_n875), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n889), .A2(new_n890), .A3(new_n861), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n920), .A2(new_n921), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n888), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n430), .B(KEYINPUT57), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n625), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n909), .A2(new_n744), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n918), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND4_X1  g745(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n932));
  INV_X1    g746(.A(new_n575), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n918), .ZN(G60));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n893), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n590), .A2(new_n591), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n918), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n940), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n923), .A2(new_n926), .A3(new_n942), .A4(new_n938), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n941), .A2(new_n943), .ZN(G63));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n215), .A2(new_n217), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n924), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n918), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n615), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n924), .A2(new_n953), .A3(new_n949), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n945), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(KEYINPUT61), .A3(new_n951), .A4(new_n950), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G66));
  NAND2_X1  g772(.A1(new_n844), .A2(new_n855), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n210), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT122), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n210), .B1(new_n445), .B2(G224), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT123), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n911), .B1(G898), .B2(new_n210), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  NAND2_X1  g780(.A1(new_n335), .A2(new_n344), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n564), .A2(new_n566), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(new_n969));
  OAI211_X1 g783(.A(new_n747), .B(new_n652), .C1(new_n753), .C2(new_n752), .ZN(new_n970));
  INV_X1    g784(.A(new_n754), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n972), .B2(new_n868), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  INV_X1    g788(.A(new_n868), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n756), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n748), .A2(new_n375), .A3(new_n595), .A4(new_n649), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n978), .A2(new_n730), .A3(new_n733), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n770), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n210), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n210), .A2(G900), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n969), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n975), .B(KEYINPUT62), .C1(new_n676), .C2(new_n656), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n677), .B2(new_n868), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n845), .A2(new_n847), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n681), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n653), .A2(new_n375), .A3(new_n988), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n984), .A2(new_n986), .B1(new_n769), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n990), .A2(new_n756), .A3(new_n770), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n210), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n969), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n210), .B1(G227), .B2(G900), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT124), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G72));
  NOR2_X1   g810(.A1(new_n346), .A2(new_n324), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI211_X1 g813(.A(KEYINPUT127), .B(new_n999), .C1(new_n980), .C2(new_n959), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n844), .A2(new_n855), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1002), .A2(new_n770), .A3(new_n979), .A4(new_n977), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT127), .B1(new_n1003), .B2(new_n999), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n997), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n951), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n346), .A2(new_n324), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1002), .A2(new_n990), .A3(new_n756), .A4(new_n770), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n999), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n877), .A2(new_n884), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1007), .A2(new_n999), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1012), .A2(new_n997), .A3(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1006), .A2(new_n1011), .A3(new_n1014), .ZN(G57));
endmodule


