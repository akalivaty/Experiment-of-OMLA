//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT67), .B1(new_n189), .B2(G116), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(new_n187), .A3(G119), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n200), .A2(KEYINPUT65), .A3(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT65), .B1(new_n200), .B2(G146), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n197), .B(new_n199), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(G143), .B2(new_n196), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n207), .B2(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  XNOR2_X1  g024(.A(G134), .B(G137), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G134), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT66), .B(G131), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n214), .B2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(KEYINPUT11), .A3(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n214), .A2(G137), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n212), .A4(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n224), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n200), .A2(G146), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n196), .B2(G143), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n200), .A2(KEYINPUT65), .A3(G146), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n197), .B2(new_n204), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT0), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n198), .A3(KEYINPUT64), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n225), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n225), .B2(new_n242), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT68), .B(new_n195), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n195), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n225), .A2(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT30), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n225), .A2(new_n242), .A3(new_n243), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n225), .A3(new_n242), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n246), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n257), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n264));
  INV_X1    g078(.A(new_n252), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n247), .B1(new_n242), .B2(new_n225), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT28), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n263), .B(new_n264), .C1(new_n262), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G902), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(KEYINPUT28), .C1(new_n265), .C2(new_n266), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n262), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n269), .B(KEYINPUT72), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n276), .A2(KEYINPUT29), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n272), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G472), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n255), .A2(new_n277), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(KEYINPUT31), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n255), .A2(new_n288), .A3(new_n277), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n270), .A2(new_n262), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(G472), .A2(G902), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n294), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT32), .B(new_n296), .C1(new_n287), .C2(new_n292), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n281), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G125), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G140), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT16), .ZN(new_n303));
  OR3_X1    g117(.A1(new_n301), .A2(KEYINPUT16), .A3(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n196), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n304), .A3(G146), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n189), .A2(G128), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n189), .A2(G128), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(KEYINPUT23), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n198), .A2(G119), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT24), .B(G110), .Z(new_n315));
  AOI22_X1  g129(.A1(new_n312), .A2(G110), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n312), .A2(G110), .B1(new_n314), .B2(new_n315), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n300), .A2(new_n302), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n307), .C1(G146), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G137), .ZN(new_n322));
  INV_X1    g136(.A(G953), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G221), .A3(G234), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n321), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n272), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G217), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(G234), .B2(new_n272), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n326), .B(new_n272), .C1(new_n330), .C2(G234), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n298), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  AOI22_X1  g154(.A1(KEYINPUT73), .A2(new_n339), .B1(new_n340), .B2(G107), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  INV_X1    g156(.A(G107), .ZN(new_n343));
  AND4_X1   g157(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT3), .A4(G104), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n342), .A2(KEYINPUT3), .B1(new_n343), .B2(G104), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n338), .B(new_n341), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n347));
  OAI22_X1  g161(.A1(KEYINPUT73), .A2(new_n339), .B1(new_n340), .B2(G107), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT3), .A4(G104), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n338), .B1(new_n350), .B2(new_n341), .ZN(new_n351));
  MUX2_X1   g165(.A(new_n347), .B(KEYINPUT4), .S(new_n351), .Z(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n241), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n340), .A2(G107), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n343), .A2(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n346), .B2(new_n357), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT10), .B(new_n209), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n346), .A2(new_n357), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n207), .A2(new_n198), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n203), .B1(new_n233), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n353), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n228), .ZN(new_n370));
  INV_X1    g184(.A(new_n228), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n353), .A2(new_n371), .A3(new_n361), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G110), .B(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n323), .A2(G227), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n374), .B(new_n375), .Z(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n378));
  INV_X1    g192(.A(new_n209), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n358), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n366), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n228), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n371), .B1(new_n380), .B2(new_n366), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(KEYINPUT12), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n376), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n385), .A3(new_n383), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n372), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(G902), .B1(new_n377), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G469), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n370), .A2(new_n372), .A3(new_n389), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n372), .A3(new_n390), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n376), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G469), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n393), .A2(new_n272), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  OAI21_X1  g216(.A(G221), .B1(new_n402), .B2(G902), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n200), .A2(KEYINPUT82), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(G214), .A3(new_n258), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(G143), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n408), .A2(new_n323), .A3(G214), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT18), .A3(G131), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n319), .B(G146), .ZN(new_n412));
  AND2_X1   g226(.A1(KEYINPUT18), .A2(G131), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n411), .B(new_n412), .C1(new_n410), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n410), .B(new_n212), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G143), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n419), .A2(new_n405), .B1(new_n258), .B2(G214), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n323), .A3(G214), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n418), .A2(G143), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT17), .B(G131), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n410), .A2(KEYINPUT85), .A3(KEYINPUT17), .A4(G131), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n308), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n417), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g244(.A(KEYINPUT86), .B(new_n308), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n414), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n340), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n414), .C1(new_n430), .C2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n272), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G475), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT19), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT19), .B1(new_n300), .B2(new_n302), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n441), .B(new_n196), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n307), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n319), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT19), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n441), .B1(new_n449), .B2(new_n196), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT84), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n415), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n196), .B1(new_n442), .B2(new_n443), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n307), .A4(new_n444), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n414), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n435), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n437), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n460), .A2(KEYINPUT87), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n459), .B2(new_n437), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT87), .B1(new_n465), .B2(new_n461), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n440), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n187), .A2(G122), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n343), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n187), .A2(G122), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(new_n476), .C1(new_n470), .C2(KEYINPUT14), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(G116), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n472), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(new_n476), .B2(KEYINPUT14), .ZN(new_n481));
  OAI211_X1 g295(.A(G107), .B(new_n477), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n198), .A2(G143), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n198), .A2(G143), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n485), .A2(G134), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n483), .B(KEYINPUT88), .ZN(new_n488));
  INV_X1    g302(.A(new_n486), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n214), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n474), .B(new_n482), .C1(new_n487), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n486), .B(KEYINPUT13), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n492), .B2(new_n485), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n473), .B(new_n343), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n214), .A3(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n402), .A2(new_n330), .A3(G953), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n491), .A2(new_n496), .A3(new_n498), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n498), .B1(new_n491), .B2(new_n496), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT90), .B(new_n272), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n203), .A2(new_n208), .A3(new_n301), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n241), .B2(new_n301), .ZN(new_n514));
  INV_X1    g328(.A(G224), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G953), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n514), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g332(.A(G113), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n188), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n518), .A2(new_n521), .B1(new_n193), .B2(new_n194), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n359), .B2(new_n360), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n351), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n195), .B(new_n525), .C1(new_n351), .C2(new_n347), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n526), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(KEYINPUT78), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n528), .A2(KEYINPUT6), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n529), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(new_n515), .B2(G953), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n514), .B(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n193), .A2(new_n194), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n359), .B2(new_n360), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT79), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n193), .A2(new_n540), .A3(KEYINPUT5), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n521), .A2(KEYINPUT80), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n521), .A2(KEYINPUT80), .ZN(new_n544));
  AND4_X1   g358(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n539), .A2(new_n545), .B1(new_n363), .B2(new_n522), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n527), .B(KEYINPUT8), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n537), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n533), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G210), .B1(G237), .B2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n533), .A2(new_n550), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G214), .B1(G237), .B2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n323), .A2(G952), .ZN(new_n560));
  NAND2_X1  g374(.A1(G234), .A2(G237), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(G902), .A3(G953), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n556), .A2(new_n559), .A3(new_n568), .ZN(new_n569));
  NOR4_X1   g383(.A1(new_n404), .A2(new_n469), .A3(new_n512), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n337), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  INV_X1    g386(.A(new_n335), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n293), .A2(new_n294), .ZN(new_n574));
  INV_X1    g388(.A(G472), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n287), .B2(new_n292), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n573), .A2(new_n404), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(KEYINPUT91), .Z(new_n579));
  OAI21_X1  g393(.A(KEYINPUT33), .B1(new_n498), .B2(KEYINPUT93), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n507), .B2(new_n508), .ZN(new_n581));
  INV_X1    g395(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n500), .A2(new_n501), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n504), .A2(G902), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n581), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n502), .B2(G478), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT95), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n469), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n554), .A2(KEYINPUT92), .A3(new_n555), .ZN(new_n595));
  INV_X1    g409(.A(new_n557), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n552), .B1(new_n533), .B2(new_n550), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n568), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n579), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  NAND2_X1  g418(.A1(new_n460), .A2(new_n462), .ZN(new_n605));
  INV_X1    g419(.A(new_n466), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n465), .A2(new_n466), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(new_n512), .A3(new_n440), .A4(new_n568), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT96), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n595), .A2(new_n599), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n607), .A2(new_n608), .B1(new_n439), .B2(G475), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n512), .A4(new_n568), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n611), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n579), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  XOR2_X1   g435(.A(new_n321), .B(KEYINPUT98), .Z(new_n622));
  INV_X1    g436(.A(KEYINPUT36), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n325), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n625), .A2(G902), .A3(new_n331), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n332), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n577), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n570), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT37), .B(G110), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G12));
  NAND2_X1  g446(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n293), .A2(new_n282), .A3(new_n294), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n404), .B1(new_n635), .B2(new_n281), .ZN(new_n636));
  INV_X1    g450(.A(new_n627), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n562), .B1(G900), .B2(new_n564), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n614), .A2(new_n512), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n612), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n636), .A2(KEYINPUT100), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n403), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n399), .B1(new_n392), .B2(new_n393), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n398), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n298), .A2(new_n644), .A3(new_n637), .A4(new_n640), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND4_X1  g463(.A1(new_n627), .A2(new_n469), .A3(new_n512), .A4(new_n557), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT101), .Z(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n638), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT70), .B1(new_n255), .B2(new_n277), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n660), .B2(G902), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n295), .B2(new_n297), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n556), .B(KEYINPUT38), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n651), .A2(new_n655), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND3_X1  g481(.A1(new_n469), .A2(new_n593), .A3(new_n638), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(KEYINPUT103), .A3(new_n613), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n668), .B2(new_n612), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n636), .A2(new_n670), .A3(new_n637), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NOR2_X1   g488(.A1(new_n392), .A2(new_n393), .ZN(new_n675));
  AOI211_X1 g489(.A(G469), .B(G902), .C1(new_n377), .C2(new_n391), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n675), .A2(new_n676), .A3(new_n642), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n298), .A2(new_n601), .A3(new_n335), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NAND4_X1  g494(.A1(new_n617), .A2(new_n298), .A3(new_n335), .A4(new_n677), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(G116), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G18));
  NOR2_X1   g497(.A1(new_n627), .A2(new_n567), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n298), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n469), .A2(new_n512), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n377), .A2(new_n391), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n272), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n403), .A3(new_n394), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n612), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n685), .A2(KEYINPUT105), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n298), .A3(new_n686), .A4(new_n684), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n291), .B1(new_n658), .B2(KEYINPUT31), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n698), .B(G472), .C1(new_n699), .C2(G902), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT107), .B1(new_n576), .B2(new_n575), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n276), .A2(new_n278), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n262), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n287), .A2(new_n704), .A3(KEYINPUT106), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n289), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT106), .B1(new_n287), .B2(new_n704), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n294), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n335), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT108), .B1(new_n469), .B2(new_n512), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n469), .A2(KEYINPUT108), .A3(new_n512), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n677), .A2(new_n568), .A3(new_n613), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n709), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n471), .ZN(G24));
  INV_X1    g530(.A(new_n707), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n289), .A3(new_n705), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n718), .A2(new_n294), .B1(new_n700), .B2(new_n701), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n637), .A3(new_n669), .A4(new_n691), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT109), .B(G125), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G27));
  AND2_X1   g536(.A1(new_n384), .A2(new_n387), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n390), .A2(new_n372), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n376), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(G469), .B(new_n727), .C1(new_n397), .C2(new_n726), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n642), .B1(new_n728), .B2(new_n643), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT111), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n556), .A2(new_n596), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n298), .A2(new_n335), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n733), .A3(new_n669), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n736), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n730), .A2(new_n733), .A3(new_n669), .A4(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n212), .ZN(G33));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n729), .B(new_n742), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n743), .A2(new_n639), .A3(new_n732), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n214), .ZN(G36));
  NOR2_X1   g559(.A1(new_n397), .A2(KEYINPUT45), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n393), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT45), .B(new_n727), .C1(new_n397), .C2(new_n726), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n400), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n394), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n750), .A2(new_n751), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n403), .B(new_n653), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  INV_X1    g571(.A(new_n469), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n593), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT43), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n577), .A2(new_n637), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n759), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n577), .A4(new_n637), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n765), .A3(new_n731), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n756), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(G137), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G39));
  OAI21_X1  g586(.A(new_n403), .B1(new_n753), .B2(new_n754), .ZN(new_n773));
  NOR2_X1   g587(.A1(KEYINPUT115), .A2(KEYINPUT47), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  OAI221_X1 g592(.A(new_n403), .B1(new_n775), .B2(new_n776), .C1(new_n753), .C2(new_n754), .ZN(new_n779));
  INV_X1    g593(.A(new_n731), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n298), .A2(new_n335), .A3(new_n668), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NOR4_X1   g597(.A1(new_n573), .A2(new_n663), .A3(new_n642), .A4(new_n558), .ZN(new_n784));
  INV_X1    g598(.A(new_n662), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n675), .A2(new_n676), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n759), .B1(new_n787), .B2(KEYINPUT49), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n760), .A2(new_n709), .A3(new_n562), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n663), .A2(new_n690), .A3(new_n557), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT122), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT50), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n690), .A2(new_n780), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n785), .A2(new_n797), .A3(new_n335), .A4(new_n563), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT123), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n799), .A2(new_n469), .A3(new_n593), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n760), .A2(new_n562), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n637), .A3(new_n719), .A4(new_n797), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n796), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n791), .A2(new_n731), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n787), .A2(new_n403), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n778), .B2(new_n779), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n778), .A2(new_n779), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n807), .B(KEYINPUT121), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n804), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n801), .A2(new_n337), .A3(new_n797), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT48), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n791), .A2(new_n691), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n560), .B(new_n816), .C1(new_n799), .C2(new_n594), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n809), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n645), .A2(new_n646), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n645), .A2(new_n646), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n673), .B(new_n720), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n638), .B(KEYINPUT119), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n627), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n662), .A2(new_n826), .A3(new_n729), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n711), .A2(new_n613), .A3(new_n712), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n825), .B1(new_n635), .B2(new_n661), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n469), .A2(KEYINPUT108), .A3(new_n512), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n710), .A3(new_n612), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .A4(new_n729), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n744), .B1(new_n737), .B2(new_n739), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n719), .A2(new_n637), .A3(new_n669), .A4(new_n731), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n743), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n637), .A2(new_n702), .A3(new_n669), .A4(new_n708), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n730), .A3(KEYINPUT118), .A4(new_n731), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n637), .A2(new_n638), .ZN(new_n843));
  INV_X1    g657(.A(new_n614), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n843), .A2(new_n512), .A3(new_n844), .A4(new_n780), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n840), .A2(new_n842), .B1(new_n636), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n836), .A2(new_n837), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n570), .B1(new_n337), .B2(new_n628), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n758), .A2(new_n512), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n569), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT117), .B1(new_n849), .B2(new_n569), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n578), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n594), .A2(new_n569), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n578), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n298), .A2(new_n335), .A3(new_n677), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n611), .A2(new_n613), .A3(new_n616), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n678), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n715), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT116), .B1(new_n859), .B2(new_n696), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(KEYINPUT116), .A3(new_n696), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n855), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n641), .A2(new_n647), .B1(new_n841), .B2(new_n691), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n829), .A2(new_n834), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n673), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n847), .A2(new_n863), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n836), .A2(new_n867), .A3(new_n837), .A4(new_n846), .ZN(new_n871));
  INV_X1    g685(.A(new_n855), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n693), .B(KEYINPUT105), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n690), .A2(new_n567), .A3(new_n612), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n335), .A3(new_n708), .A4(new_n702), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n681), .B(new_n678), .C1(new_n875), .C2(new_n713), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n872), .B1(new_n878), .B2(new_n860), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n868), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n820), .B1(new_n870), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n837), .A2(new_n846), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n864), .A2(new_n865), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n859), .A2(new_n696), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n848), .A2(new_n852), .A3(KEYINPUT53), .A4(new_n854), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n882), .A2(new_n886), .A3(new_n867), .A4(new_n836), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n880), .A2(new_n820), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n819), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n790), .B1(new_n889), .B2(new_n890), .ZN(G75));
  AOI21_X1  g705(.A(new_n272), .B1(new_n880), .B2(new_n887), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G210), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n531), .A2(new_n532), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n517), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n323), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n895), .A2(new_n898), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(G51));
  AOI21_X1  g718(.A(new_n820), .B1(new_n880), .B2(new_n887), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n888), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n399), .B(KEYINPUT57), .Z(new_n907));
  OAI21_X1  g721(.A(new_n687), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n892), .A2(new_n748), .A3(new_n747), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n892), .A2(new_n460), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n460), .B1(new_n892), .B2(new_n911), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n914), .A2(new_n915), .A3(new_n900), .A4(new_n916), .ZN(G60));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n581), .A2(new_n583), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n880), .A2(new_n887), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n880), .A2(new_n887), .A3(new_n820), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n918), .B1(new_n925), .B2(new_n900), .ZN(new_n926));
  OAI211_X1 g740(.A(KEYINPUT125), .B(new_n901), .C1(new_n906), .C2(new_n921), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n920), .B1(new_n881), .B2(new_n888), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n581), .A2(new_n583), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n927), .A3(new_n930), .ZN(G63));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n326), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n900), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n625), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n937), .B(KEYINPUT61), .C1(new_n625), .C2(new_n935), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n566), .B2(new_n515), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n863), .B2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n896), .B1(G898), .B2(new_n323), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G69));
  NOR2_X1   g760(.A1(new_n244), .A2(new_n245), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(new_n449), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n782), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n770), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n756), .A2(new_n337), .A3(new_n832), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n837), .ZN(new_n953));
  INV_X1    g767(.A(new_n823), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n323), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(G900), .A2(G953), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n654), .B1(new_n594), .B2(new_n849), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n733), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n782), .B(new_n959), .C1(new_n768), .C2(new_n769), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n954), .A2(new_n666), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n964), .A2(G953), .A3(new_n948), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n323), .B1(G227), .B2(G900), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(new_n870), .A2(new_n880), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n575), .A2(new_n272), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n658), .B2(new_n263), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n256), .A2(new_n277), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n964), .A2(new_n863), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n976), .B(new_n978), .C1(new_n979), .C2(new_n973), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n951), .A2(new_n954), .A3(new_n953), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n981), .B2(new_n879), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n256), .A2(new_n277), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n900), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n973), .B1(new_n964), .B2(new_n863), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT127), .B1(new_n985), .B2(new_n977), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n975), .A2(new_n980), .A3(new_n984), .A4(new_n986), .ZN(G57));
endmodule


