//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n462), .A2(G136), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n459), .B2(new_n460), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n482), .B(new_n485), .C1(new_n460), .C2(new_n459), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(G126), .B2(new_n475), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  NAND2_X1  g068(.A1(KEYINPUT67), .A2(G543), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n501), .A2(new_n507), .ZN(G166));
  INV_X1    g083(.A(new_n503), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G89), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n498), .A2(G63), .A3(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(G51), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n511), .B(new_n513), .C1(new_n505), .C2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(G168));
  AOI22_X1  g091(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(new_n500), .ZN(new_n518));
  INV_X1    g093(.A(G90), .ZN(new_n519));
  INV_X1    g094(.A(G52), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n503), .A2(new_n519), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G171));
  NAND3_X1  g097(.A1(new_n498), .A2(new_n502), .A3(G81), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT68), .B(G43), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n502), .A2(new_n524), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n523), .B2(new_n525), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n500), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G860), .A3(new_n532), .ZN(G153));
  NAND4_X1  g108(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g109(.A1(G1), .A2(G3), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT8), .ZN(new_n536));
  NAND4_X1  g111(.A1(G319), .A2(G483), .A3(G661), .A4(new_n536), .ZN(G188));
  INV_X1    g112(.A(G53), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n505), .A2(KEYINPUT9), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT9), .B1(new_n505), .B2(new_n538), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(new_n540), .B1(G91), .B2(new_n509), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n498), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n500), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n545));
  NOR3_X1   g120(.A1(new_n542), .A2(new_n545), .A3(new_n500), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n541), .B(KEYINPUT71), .C1(new_n544), .C2(new_n546), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G299));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g128(.A1(G171), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n518), .B2(new_n521), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  NAND2_X1  g134(.A1(new_n509), .A2(G87), .ZN(new_n560));
  INV_X1    g135(.A(new_n505), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G49), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(G288));
  NAND2_X1  g139(.A1(new_n498), .A2(G61), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n500), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n509), .A2(G86), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  AOI22_X1  g146(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n500), .ZN(new_n573));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n503), .A2(new_n574), .B1(new_n505), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(new_n509), .A2(G92), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT10), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(G54), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n498), .A2(G66), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT74), .Z(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  MUX2_X1   g166(.A(G301), .B(new_n590), .S(new_n591), .Z(G284));
  MUX2_X1   g167(.A(G301), .B(new_n590), .S(new_n591), .Z(G321));
  NOR2_X1   g168(.A1(G286), .A2(new_n591), .ZN(new_n594));
  XOR2_X1   g169(.A(G299), .B(KEYINPUT75), .Z(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n591), .ZN(G297));
  AOI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(new_n591), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G860), .ZN(G148));
  OAI21_X1  g174(.A(new_n532), .B1(new_n527), .B2(new_n529), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n590), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n591), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g179(.A(KEYINPUT3), .B(G2104), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n464), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(G2100), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n462), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n475), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n463), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2430), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n623), .A2(KEYINPUT76), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(KEYINPUT76), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n624), .A2(new_n625), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n632), .ZN(new_n634));
  AND3_X1   g209(.A1(new_n633), .A2(new_n634), .A3(G14), .ZN(G401));
  XNOR2_X1  g210(.A(G2084), .B(G2090), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT77), .Z(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n638), .B(KEYINPUT17), .Z(new_n641));
  INV_X1    g216(.A(new_n639), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n636), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n636), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n639), .A2(new_n636), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n659), .B(new_n661), .C1(new_n654), .C2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XOR2_X1   g238(.A(G1981), .B(G1986), .Z(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT78), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n663), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G4), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n589), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1348), .ZN(new_n674));
  NOR2_X1   g249(.A1(G168), .A2(new_n671), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(G21), .ZN(new_n676));
  INV_X1    g251(.A(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(G171), .A2(new_n671), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(G5), .B2(new_n671), .ZN(new_n679));
  INV_X1    g254(.A(G1961), .ZN(new_n680));
  AOI22_X1  g255(.A1(new_n676), .A2(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(G19), .B(new_n600), .S(G16), .Z(new_n682));
  OAI221_X1 g257(.A(new_n681), .B1(new_n680), .B2(new_n679), .C1(new_n682), .C2(G1341), .ZN(new_n683));
  AOI211_X1 g258(.A(new_n674), .B(new_n683), .C1(G1341), .C2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(G299), .A2(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n671), .A2(G20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT23), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1956), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n475), .A2(G129), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n464), .A2(G105), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G141), .B2(new_n462), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT26), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n700), .B2(G32), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(G33), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT25), .Z(new_n710));
  INV_X1    g285(.A(new_n462), .ZN(new_n711));
  INV_X1    g286(.A(G139), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT88), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n605), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n463), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(new_n700), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G2072), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n700), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n700), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n707), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G11), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT30), .B(G28), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n700), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n700), .B2(new_n616), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  INV_X1    g306(.A(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n732), .B2(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(KEYINPUT24), .B2(new_n732), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n470), .B2(new_n700), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n730), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n702), .B2(new_n704), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n700), .A2(G35), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n700), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2090), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n731), .B2(new_n735), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n718), .A2(G2072), .B1(new_n723), .B2(new_n722), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n705), .A2(new_n706), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n700), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n462), .A2(G140), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G116), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G128), .B2(new_n475), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n700), .ZN(new_n759));
  INV_X1    g334(.A(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT92), .B1(new_n676), .B2(new_n677), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n676), .A2(KEYINPUT92), .A3(new_n677), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n748), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n747), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n684), .A2(new_n690), .A3(new_n725), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n671), .A2(G22), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT84), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G166), .B2(new_n671), .ZN(new_n770));
  INV_X1    g345(.A(G1971), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(KEYINPUT85), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(KEYINPUT85), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G23), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT83), .Z(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G288), .B2(new_n671), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT33), .B(G1976), .Z(new_n778));
  XOR2_X1   g353(.A(new_n777), .B(new_n778), .Z(new_n779));
  NOR3_X1   g354(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n671), .A2(G6), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G305), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT82), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n671), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n577), .B2(new_n671), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  AND3_X1   g368(.A1(new_n700), .A2(KEYINPUT80), .A3(G25), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT80), .B1(new_n700), .B2(G25), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n462), .A2(G131), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n475), .A2(G119), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n463), .A2(G107), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n796), .B(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n794), .B(new_n795), .C1(new_n804), .C2(G29), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n792), .B1(new_n793), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n793), .B2(new_n805), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n787), .A2(new_n788), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n766), .B1(new_n767), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n767), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n810), .B1(new_n809), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(G311));
  AND3_X1   g389(.A1(new_n809), .A2(KEYINPUT98), .A3(new_n811), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT98), .B1(new_n809), .B2(new_n811), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n589), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT38), .Z(new_n820));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n530), .A2(new_n821), .A3(new_n532), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n600), .A2(KEYINPUT99), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n500), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n503), .A2(new_n827), .B1(new_n505), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n822), .A2(new_n823), .A3(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n820), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n818), .B1(new_n836), .B2(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT100), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n840), .A3(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n831), .A2(G860), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT101), .ZN(G145));
  XNOR2_X1  g421(.A(new_n616), .B(new_n470), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n479), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n475), .A2(G126), .ZN(new_n850));
  INV_X1    g425(.A(new_n490), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n486), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n485), .B1(new_n605), .B2(new_n482), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT102), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n484), .A2(new_n856), .A3(new_n486), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n852), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n758), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n717), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n484), .A2(new_n856), .A3(new_n486), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n484), .B2(new_n486), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n491), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n758), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n717), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n698), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n860), .A2(new_n866), .A3(new_n699), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n475), .A2(G130), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n463), .A2(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G142), .B2(new_n462), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n607), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(new_n804), .Z(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n868), .A2(new_n877), .A3(new_n869), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n849), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n868), .A2(KEYINPUT104), .A3(new_n877), .A4(new_n869), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n848), .B(KEYINPUT105), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n885), .A2(new_n879), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n883), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G395));
  XNOR2_X1  g469(.A(new_n834), .B(new_n602), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n590), .B1(new_n549), .B2(new_n551), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n547), .A2(new_n548), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n550), .A3(new_n589), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(new_n577), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(G288), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(KEYINPUT42), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n902), .B(new_n904), .C1(new_n911), .C2(KEYINPUT42), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n907), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n907), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n830), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n830), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n556), .A2(G168), .ZN(new_n921));
  OR2_X1    g496(.A1(G168), .A2(G171), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n832), .A2(new_n833), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n903), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n833), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n830), .B1(new_n822), .B2(new_n823), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n921), .B(new_n922), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n832), .B2(new_n833), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n924), .ZN(new_n934));
  OAI22_X1  g509(.A1(new_n899), .A2(new_n900), .B1(new_n934), .B2(new_n930), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n935), .A3(new_n910), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n889), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  INV_X1    g513(.A(new_n910), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n929), .A2(new_n932), .A3(new_n924), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT41), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n903), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n899), .A2(KEYINPUT108), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n925), .A2(new_n928), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n910), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n936), .A2(new_n889), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT43), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n919), .B1(new_n941), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n937), .B2(new_n940), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n939), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n937), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n951), .B2(new_n952), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n954), .B1(new_n962), .B2(new_n919), .ZN(G397));
  XNOR2_X1  g538(.A(new_n758), .B(new_n760), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(G1996), .B2(new_n698), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n863), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n465), .A2(G40), .A3(new_n469), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT112), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n699), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n804), .B(new_n793), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n971), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n577), .A2(new_n791), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT111), .Z(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n791), .B2(new_n577), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT50), .B1(new_n858), .B2(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n487), .B2(new_n491), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n985), .A2(KEYINPUT119), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT119), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n984), .B(new_n970), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n689), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n863), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n853), .A2(new_n854), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n852), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n969), .B1(new_n994), .B2(new_n968), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT56), .B(G2072), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n991), .A2(new_n995), .A3(KEYINPUT122), .A4(new_n996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n990), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n547), .B(KEYINPUT57), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n855), .A2(new_n857), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n1004), .B2(new_n491), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n760), .A3(new_n970), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n863), .A2(new_n986), .A3(new_n992), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n863), .A2(new_n1008), .A3(new_n986), .A4(new_n992), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n969), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(G1348), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT123), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n589), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1013), .B2(new_n589), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1003), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT124), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1021), .B(new_n1003), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT60), .B(new_n1006), .C1(new_n1012), .C2(G1348), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT125), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n589), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1026), .A3(new_n590), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT61), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1003), .A2(KEYINPUT61), .A3(new_n1016), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n991), .A2(new_n995), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n1038), .A2(G1996), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1005), .A2(new_n970), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT58), .B(G1341), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n600), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1036), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1020), .B(new_n1022), .C1(new_n1032), .C2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G288), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G1976), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1040), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1050), .A2(G1976), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1052), .A2(KEYINPUT52), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n568), .A2(new_n569), .A3(new_n1055), .A4(new_n570), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(G86), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n503), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n570), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n567), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1056), .B(KEYINPUT49), .C1(new_n1060), .C2(new_n1055), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1061), .A2(new_n1040), .A3(new_n1049), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1056), .B1(new_n1060), .B2(new_n1055), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1062), .A2(new_n1065), .B1(new_n1052), .B2(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n863), .A2(new_n992), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n969), .B1(new_n1067), .B2(KEYINPUT50), .ZN(new_n1068));
  INV_X1    g643(.A(G2090), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1068), .B(new_n1069), .C1(new_n988), .C2(new_n987), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1038), .A2(new_n771), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1048), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G166), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT55), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1054), .B(new_n1066), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n969), .A2(G2090), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(KEYINPUT114), .B(new_n1078), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1082));
  OAI211_X1 g657(.A(G8), .B(new_n1075), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT113), .B1(new_n985), .B2(new_n986), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n986), .B2(new_n1005), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1011), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1077), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n1071), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(G8), .A4(new_n1075), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1076), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1038), .B2(G2078), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1012), .B2(G1961), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT45), .B1(new_n863), .B2(new_n992), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n1098), .B2(new_n969), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n970), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1095), .A2(G2078), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n556), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n970), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n680), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1103), .B1(new_n969), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1108), .B2(new_n969), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n967), .A2(new_n968), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n991), .A3(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1107), .A2(G301), .A3(new_n1096), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1107), .A2(G301), .A3(new_n1096), .A4(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1112), .B(new_n1096), .C1(new_n1012), .C2(G1961), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1118), .B2(G171), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1114), .A2(new_n1115), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G168), .A2(new_n1048), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1123), .A2(new_n677), .B1(new_n1012), .B2(new_n731), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1122), .B1(new_n1124), .B2(new_n1073), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n677), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1012), .A2(new_n731), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1049), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1125), .B(KEYINPUT51), .C1(new_n1129), .C2(G168), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1131), .A3(new_n1122), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1094), .A2(new_n1120), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1047), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1130), .A2(KEYINPUT62), .A3(new_n1132), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1105), .B(new_n1076), .C1(new_n1084), .C2(new_n1093), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1084), .A2(new_n1093), .A3(new_n1054), .A4(new_n1066), .ZN(new_n1141));
  AOI211_X1 g716(.A(G1976), .B(G288), .C1(new_n1062), .C2(new_n1065), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1056), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1049), .B(new_n1040), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT118), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1141), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1134), .A2(new_n1140), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1128), .A2(G168), .A3(new_n1049), .ZN(new_n1152));
  AOI211_X1 g727(.A(new_n1076), .B(new_n1152), .C1(new_n1084), .C2(new_n1093), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1153), .B2(KEYINPUT63), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1152), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1094), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(KEYINPUT121), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1075), .B1(new_n1091), .B2(G8), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1066), .A2(new_n1054), .ZN(new_n1160));
  NOR4_X1   g735(.A1(new_n1159), .A2(new_n1152), .A3(new_n1157), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1154), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n983), .B1(new_n1150), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n802), .A2(new_n793), .A3(new_n803), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n975), .A2(new_n1166), .B1(new_n760), .B2(new_n758), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n971), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(KEYINPUT127), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n978), .B1(new_n964), .B2(new_n698), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT46), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n974), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n974), .A2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT47), .Z(new_n1175));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1167), .A2(new_n1176), .A3(new_n971), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n980), .A2(new_n978), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT48), .Z(new_n1179));
  NOR2_X1   g754(.A1(new_n977), .A2(new_n1179), .ZN(new_n1180));
  NOR4_X1   g755(.A1(new_n1169), .A2(new_n1175), .A3(new_n1177), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g757(.A1(new_n651), .A2(G319), .ZN(new_n1184));
  NOR3_X1   g758(.A1(G401), .A2(G229), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g759(.A(new_n881), .B(KEYINPUT103), .ZN(new_n1186));
  OAI221_X1 g760(.A(new_n1185), .B1(new_n941), .B2(new_n953), .C1(new_n1186), .C2(new_n890), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


