//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  AND3_X1   g001(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  OR2_X1    g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n217), .A2(new_n219), .A3(new_n212), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n223), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n233), .A2(new_n212), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n215), .A3(new_n216), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n235), .B2(new_n236), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n234), .A2(new_n237), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n224), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n246), .B(new_n247), .C1(new_n207), .C2(new_n208), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n248), .B2(KEYINPUT28), .ZN(new_n249));
  OR2_X1    g048(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT28), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(KEYINPUT67), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n245), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n252), .A2(new_n246), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n243), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G127gat), .B(G134gat), .Z(new_n258));
  OR2_X1    g057(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G127gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT70), .A3(G134gat), .ZN(new_n265));
  OAI221_X1 g064(.A(new_n265), .B1(new_n260), .B2(KEYINPUT1), .C1(new_n258), .C2(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n257), .B(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G227gat), .A2(G233gat), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n268), .A2(KEYINPUT34), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT34), .B1(new_n268), .B2(new_n269), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n271), .A2(KEYINPUT73), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT73), .B1(new_n271), .B2(new_n272), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G71gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G99gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n268), .A2(new_n269), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n279), .B(KEYINPUT32), .C1(new_n280), .C2(new_n278), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n275), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(new_n273), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n202), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT36), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT36), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n202), .B(new_n291), .C1(new_n286), .C2(new_n288), .ZN(new_n292));
  XOR2_X1   g091(.A(G78gat), .B(G106gat), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT31), .ZN(new_n294));
  INV_X1    g093(.A(G50gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT2), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G155gat), .B(G162gat), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n304), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(KEYINPUT22), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n307), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n307), .A2(new_n319), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n315), .B1(new_n321), .B2(new_n316), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n299), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n322), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n304), .B(new_n305), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n314), .A2(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n299), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT82), .B(G22gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n323), .B2(new_n329), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n297), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n323), .B2(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT83), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n296), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n331), .B1(new_n336), .B2(KEYINPUT83), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT4), .B1(new_n267), .B2(new_n325), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n307), .A2(new_n349), .A3(new_n266), .A4(new_n263), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n321), .A2(new_n326), .A3(new_n267), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n267), .B(new_n325), .ZN(new_n357));
  INV_X1    g156(.A(new_n352), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n347), .B(new_n356), .C1(new_n360), .C2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(new_n356), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n355), .B1(new_n354), .B2(new_n359), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n346), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n232), .A2(new_n371), .A3(new_n256), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n232), .B2(new_n256), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n243), .A2(new_n249), .A3(new_n255), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n226), .A2(new_n228), .A3(new_n227), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n379), .A2(new_n212), .A3(new_n219), .A4(new_n217), .ZN(new_n380));
  AND4_X1   g179(.A1(new_n214), .A2(new_n219), .A3(new_n217), .A4(new_n220), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n380), .A2(new_n223), .B1(new_n381), .B2(new_n210), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n375), .B(KEYINPUT75), .Z(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT76), .B1(new_n378), .B2(new_n382), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n232), .A2(new_n256), .A3(new_n371), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n316), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n389), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n377), .A2(new_n315), .A3(new_n386), .A4(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n376), .A3(new_n388), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n383), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT77), .A3(new_n314), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n314), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G8gat), .B(G36gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G64gat), .ZN(new_n400));
  INV_X1    g199(.A(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n391), .A2(new_n395), .A3(new_n398), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n398), .A3(new_n395), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n402), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n404), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n369), .A2(new_n407), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n290), .A2(new_n292), .B1(new_n341), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n369), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n389), .A2(KEYINPUT78), .A3(new_n375), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT78), .B1(new_n389), .B2(new_n375), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n415), .A2(new_n416), .A3(new_n385), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT86), .B1(new_n417), .B2(new_n315), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n392), .A2(new_n393), .A3(new_n315), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n377), .A2(new_n386), .A3(new_n390), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n314), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT37), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n391), .A2(new_n425), .A3(new_n398), .A4(new_n395), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(new_n402), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT38), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n408), .A2(KEYINPUT37), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n427), .A2(KEYINPUT38), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n414), .B(new_n404), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n340), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT39), .B1(new_n357), .B2(new_n358), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT85), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n351), .A2(new_n353), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n358), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n347), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(KEYINPUT39), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(KEYINPUT40), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n361), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT40), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n409), .A3(new_n411), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n407), .A2(new_n409), .A3(KEYINPUT84), .A4(new_n411), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n440), .B(new_n442), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n413), .B1(new_n432), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n445), .A2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n287), .B1(new_n273), .B2(new_n274), .ZN(new_n450));
  INV_X1    g249(.A(new_n273), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n285), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n340), .A3(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n453), .A2(KEYINPUT35), .A3(new_n414), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT35), .B1(new_n412), .B2(new_n453), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT87), .B(KEYINPUT35), .C1(new_n412), .C2(new_n453), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n448), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n448), .B2(new_n461), .ZN(new_n464));
  NOR2_X1   g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n465), .A2(KEYINPUT14), .ZN(new_n466));
  INV_X1    g265(.A(new_n465), .ZN(new_n467));
  INV_X1    g266(.A(G29gat), .ZN(new_n468));
  INV_X1    g267(.A(G36gat), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  XOR2_X1   g271(.A(G43gat), .B(G50gat), .Z(new_n473));
  AND2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n470), .A2(new_n467), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT17), .ZN(new_n480));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT16), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(G1gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G1gat), .B2(new_n481), .ZN(new_n485));
  INV_X1    g284(.A(G8gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(KEYINPUT90), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n479), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT18), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n489), .B(new_n479), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n492), .B(KEYINPUT13), .Z(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT18), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n501));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G169gat), .B(G197gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT12), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n493), .A2(new_n506), .A3(new_n496), .A4(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n463), .A2(new_n464), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G85gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT96), .B1(new_n513), .B2(new_n401), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(G85gat), .A3(G92gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518));
  AOI22_X1  g317(.A1(KEYINPUT8), .A2(new_n518), .B1(new_n513), .B2(new_n401), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT96), .B(new_n520), .C1(new_n513), .C2(new_n401), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G99gat), .B(G106gat), .Z(new_n523));
  OR2_X1    g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n480), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n479), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT41), .ZN(new_n530));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G134gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n530), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT95), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n302), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n535), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT91), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(G71gat), .ZN(new_n544));
  INV_X1    g343(.A(G78gat), .ZN(new_n545));
  OAI221_X1 g344(.A(new_n541), .B1(new_n542), .B2(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(KEYINPUT9), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n549));
  OAI21_X1  g348(.A(G64gat), .B1(new_n549), .B2(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(KEYINPUT93), .A2(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n549), .A2(KEYINPUT93), .A3(G57gat), .A4(G64gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G127gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n489), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n557), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT94), .B(G155gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n564), .A2(new_n569), .A3(new_n565), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n539), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n512), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n524), .A3(new_n525), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT10), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT97), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n546), .A2(new_n554), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n526), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n528), .A2(new_n583), .A3(KEYINPUT10), .A4(new_n555), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT98), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n577), .A2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G176gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G204gat), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n576), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n414), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g399(.A1(new_n482), .A2(new_n486), .ZN(new_n601));
  NOR4_X1   g400(.A1(new_n576), .A2(new_n597), .A3(new_n449), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n482), .A2(new_n486), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT42), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n449), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n486), .B1(new_n598), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n603), .B2(new_n602), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n606), .B1(new_n609), .B2(new_n605), .ZN(G1325gat));
  NOR2_X1   g409(.A1(new_n286), .A2(new_n288), .ZN(new_n611));
  AOI21_X1  g410(.A(G15gat), .B1(new_n598), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n290), .A2(new_n292), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(G15gat), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n598), .B2(new_n615), .ZN(G1326gat));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n341), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT43), .B(G22gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(G1327gat));
  XNOR2_X1  g418(.A(new_n573), .B(KEYINPUT99), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n597), .B(KEYINPUT100), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n510), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT101), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n412), .A2(new_n341), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n613), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n431), .A2(new_n340), .ZN(new_n626));
  INV_X1    g425(.A(new_n440), .ZN(new_n627));
  INV_X1    g426(.A(new_n442), .ZN(new_n628));
  INV_X1    g427(.A(new_n445), .ZN(new_n629));
  INV_X1    g428(.A(new_n446), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n625), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n456), .A2(new_n457), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n633), .A2(new_n459), .B1(new_n449), .B2(new_n454), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT88), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n448), .A2(new_n461), .A3(new_n462), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n535), .B(new_n538), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT44), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n455), .B(new_n640), .C1(new_n458), .C2(new_n460), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n634), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n448), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n623), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(G29gat), .B1(new_n648), .B2(new_n369), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n636), .A3(new_n510), .A4(new_n637), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n573), .A2(new_n597), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n651), .A2(new_n369), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n654), .B2(new_n468), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n654), .A2(new_n650), .A3(new_n468), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(G1328gat));
  NOR2_X1   g456(.A1(new_n651), .A2(new_n653), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n449), .A2(G36gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n664), .B2(KEYINPUT46), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT46), .ZN(new_n666));
  OAI21_X1  g465(.A(G36gat), .B1(new_n648), .B2(new_n449), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n662), .A2(new_n668), .A3(new_n669), .A4(new_n663), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n665), .A2(new_n666), .A3(new_n667), .A4(new_n670), .ZN(G1329gat));
  INV_X1    g470(.A(G43gat), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n647), .B2(new_n614), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n658), .A2(new_n672), .A3(new_n611), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1330gat));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n512), .A2(new_n679), .A3(new_n637), .A4(new_n652), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n651), .B2(new_n653), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n680), .A2(new_n681), .A3(new_n295), .A4(new_n341), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n295), .B1(new_n647), .B2(new_n341), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT107), .B(KEYINPUT48), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n639), .A2(new_n646), .ZN(new_n686));
  INV_X1    g485(.A(new_n623), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n341), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G50gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n690));
  OR2_X1    g489(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .A4(new_n682), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n685), .A2(new_n692), .ZN(G1331gat));
  NOR2_X1   g492(.A1(new_n574), .A2(new_n510), .ZN(new_n694));
  INV_X1    g493(.A(new_n621), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT108), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n461), .A2(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n641), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n448), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n414), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT92), .B(G57gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1332gat));
  NAND2_X1  g502(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n607), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1333gat));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n544), .A3(new_n611), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n700), .A2(new_n614), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n544), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g511(.A1(new_n700), .A2(new_n341), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT110), .B(G78gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n573), .A2(new_n510), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n597), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n639), .B2(new_n646), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722), .B2(new_n369), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n539), .B1(new_n699), .B2(new_n448), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT51), .B1(new_n724), .B2(new_n716), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AND4_X1   g525(.A1(KEYINPUT51), .A2(new_n644), .A3(new_n637), .A4(new_n716), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n513), .A3(new_n597), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n723), .B1(new_n730), .B2(new_n369), .ZN(G1336gat));
  NOR2_X1   g530(.A1(new_n449), .A2(G92gat), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n695), .B(new_n732), .C1(new_n725), .C2(new_n727), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n449), .B(new_n720), .C1(new_n639), .C2(new_n646), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n401), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT52), .ZN(new_n737));
  OAI21_X1  g536(.A(G92gat), .B1(new_n722), .B2(new_n449), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n738), .A2(new_n734), .A3(new_n739), .A4(new_n733), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n722), .B2(new_n613), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n718), .A2(new_n286), .A3(G99gat), .A4(new_n288), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT112), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(G1338gat));
  INV_X1    g545(.A(G106gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n721), .B2(new_n341), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n729), .A2(new_n695), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n341), .A2(new_n747), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n621), .B(new_n752), .C1(new_n726), .C2(new_n728), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT53), .B1(new_n754), .B2(new_n748), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1339gat));
  NOR2_X1   g555(.A1(new_n491), .A2(new_n492), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n494), .A2(new_n495), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n505), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n597), .A2(new_n509), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n579), .A2(new_n582), .A3(new_n587), .A4(new_n584), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n589), .A2(KEYINPUT54), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n585), .A2(new_n763), .A3(new_n588), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n762), .A2(KEYINPUT55), .A3(new_n594), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n595), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n762), .A2(new_n594), .A3(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n510), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n637), .B1(new_n760), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n770), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n509), .A2(new_n759), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n539), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n620), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n694), .A2(new_n718), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n453), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n449), .A2(new_n414), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n510), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G113gat), .ZN(G1340gat));
  OAI21_X1  g583(.A(G120gat), .B1(new_n781), .B2(new_n621), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n718), .A2(G120gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT113), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n781), .B2(new_n787), .ZN(G1341gat));
  NOR3_X1   g587(.A1(new_n781), .A2(new_n264), .A3(new_n620), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n573), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n264), .B2(new_n790), .ZN(G1342gat));
  NAND2_X1  g590(.A1(new_n782), .A2(new_n637), .ZN(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(G1343gat));
  AOI21_X1  g595(.A(new_n340), .B1(new_n776), .B2(new_n777), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n779), .A2(new_n614), .ZN(new_n800));
  INV_X1    g599(.A(new_n573), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n768), .A2(KEYINPUT115), .A3(new_n769), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n768), .B2(new_n769), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n804), .B2(new_n766), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n767), .B(new_n806), .C1(new_n802), .C2(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n510), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n760), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n637), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n811), .B2(new_n775), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n340), .B1(new_n812), .B2(new_n777), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n799), .B(new_n800), .C1(new_n813), .C2(new_n798), .ZN(new_n814));
  OAI21_X1  g613(.A(G141gat), .B1(new_n814), .B2(new_n511), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n800), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n817), .A2(G141gat), .A3(new_n511), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n822), .A2(new_n815), .A3(new_n823), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n820), .A2(new_n821), .B1(new_n824), .B2(new_n816), .ZN(G1344gat));
  NOR2_X1   g624(.A1(new_n813), .A2(KEYINPUT57), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(G148gat), .A3(new_n597), .A4(new_n800), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n817), .A2(new_n718), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(G148gat), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n814), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT59), .B1(new_n832), .B2(new_n597), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n831), .A2(KEYINPUT59), .B1(G148gat), .B2(new_n833), .ZN(G1345gat));
  INV_X1    g633(.A(new_n817), .ZN(new_n835));
  AOI21_X1  g634(.A(G155gat), .B1(new_n835), .B2(new_n573), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n620), .A2(new_n301), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT119), .Z(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n832), .B2(new_n838), .ZN(G1346gat));
  AOI21_X1  g638(.A(G162gat), .B1(new_n835), .B2(new_n637), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n539), .A2(new_n302), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n832), .B2(new_n841), .ZN(G1347gat));
  NAND2_X1  g641(.A1(new_n607), .A2(new_n369), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n778), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n511), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n215), .ZN(G1348gat));
  NOR3_X1   g646(.A1(new_n845), .A2(new_n216), .A3(new_n621), .ZN(new_n848));
  INV_X1    g647(.A(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n597), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n216), .B2(new_n850), .ZN(G1349gat));
  OAI21_X1  g650(.A(G183gat), .B1(new_n845), .B2(new_n620), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n573), .A2(new_n246), .A3(new_n247), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g654(.A1(new_n849), .A2(new_n637), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G190gat), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT120), .A3(new_n858), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n856), .A2(G190gat), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n207), .A2(new_n208), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n859), .B(new_n862), .C1(new_n863), .C2(new_n856), .ZN(G1351gat));
  NOR2_X1   g663(.A1(new_n843), .A2(new_n614), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n797), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT121), .ZN(new_n867));
  INV_X1    g666(.A(G197gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n797), .A2(new_n869), .A3(new_n865), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(new_n868), .A3(new_n510), .A4(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n510), .B(new_n865), .C1(new_n826), .C2(new_n827), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G197gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT123), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1352gat));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n828), .A2(new_n865), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n621), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n828), .A2(KEYINPUT124), .A3(new_n695), .A4(new_n865), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(G204gat), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n866), .A2(G204gat), .A3(new_n718), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT62), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1353gat));
  OAI21_X1  g687(.A(G211gat), .B1(new_n882), .B2(new_n801), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT63), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(G211gat), .C1(new_n882), .C2(new_n801), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n309), .A3(new_n573), .A4(new_n870), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT125), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(G1354gat));
  NOR3_X1   g694(.A1(new_n882), .A2(new_n310), .A3(new_n539), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n867), .A2(new_n637), .A3(new_n870), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(new_n310), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(KEYINPUT126), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(KEYINPUT126), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(G1355gat));
endmodule


