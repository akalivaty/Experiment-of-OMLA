//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(new_n206), .A2(G50), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n212), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n229));
  AND3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n213), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n223), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n218), .B(new_n232), .C1(new_n224), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G179), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT70), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  INV_X1    g0064(.A(new_n221), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n257), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(G1698), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n276), .B1(new_n277), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n270), .A2(new_n283), .A3(KEYINPUT71), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT71), .B1(new_n270), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n251), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n270), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n270), .A2(new_n283), .A3(KEYINPUT71), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n293));
  INV_X1    g0093(.A(G150), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n212), .A2(G33), .ZN(new_n297));
  XOR2_X1   g0097(.A(KEYINPUT8), .B(G58), .Z(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n293), .B1(new_n294), .B2(new_n296), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n221), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(new_n211), .B2(G20), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(G50), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n286), .A2(new_n292), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT9), .B1(new_n303), .B2(new_n307), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  INV_X1    g0112(.A(new_n307), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n300), .C2(new_n302), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n289), .A2(G200), .A3(new_n291), .ZN(new_n316));
  OAI21_X1  g0116(.A(G190), .B1(new_n284), .B2(new_n285), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n317), .A3(new_n316), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT10), .A3(new_n319), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n310), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n214), .A2(G1), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n212), .A2(G68), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT73), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n306), .A2(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT74), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n326), .B1(G50), .B2(new_n295), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n277), .B2(new_n297), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n302), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT11), .Z(new_n335));
  NOR2_X1   g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n256), .A2(G238), .A3(new_n260), .A4(new_n258), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n269), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n275), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n338), .B(new_n341), .C1(new_n344), .C2(new_n258), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n258), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n290), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n347), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n251), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n348), .A2(new_n349), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n337), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(G200), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n336), .B(new_n354), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n261), .A2(G244), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n358), .A2(new_n269), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n278), .A2(G232), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G107), .ZN(new_n362));
  INV_X1    g0162(.A(G238), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n361), .B1(new_n362), .B2(new_n278), .C1(new_n280), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n282), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n359), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n251), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n306), .A2(G77), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(G77), .B2(new_n304), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G20), .A2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n297), .B2(new_n372), .C1(new_n299), .C2(new_n296), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n302), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n366), .B2(new_n290), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n366), .A2(G200), .ZN(new_n378));
  INV_X1    g0178(.A(new_n374), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n367), .B2(G190), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n324), .A2(new_n357), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n304), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n298), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n306), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n298), .ZN(new_n386));
  INV_X1    g0186(.A(new_n302), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n204), .A2(new_n205), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n202), .A2(new_n203), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n295), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(KEYINPUT3), .A2(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n212), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n274), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n273), .A2(new_n212), .A3(new_n274), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n203), .B1(new_n404), .B2(new_n397), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n392), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n387), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n397), .A2(KEYINPUT76), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n395), .A2(new_n410), .A3(KEYINPUT7), .A4(new_n212), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n411), .A3(new_n404), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  INV_X1    g0213(.A(new_n392), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n386), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n256), .A2(G232), .A3(new_n260), .A4(new_n258), .ZN(new_n419));
  MUX2_X1   g0219(.A(G223), .B(G226), .S(G1698), .Z(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n278), .B1(G33), .B2(G87), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n269), .C1(new_n421), .C2(new_n258), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n251), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(G169), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT18), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G200), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G190), .B2(new_n422), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n405), .A2(KEYINPUT75), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n400), .B(new_n203), .C1(new_n404), .C2(new_n397), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT16), .B(new_n414), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n417), .A2(new_n432), .A3(new_n302), .ZN(new_n433));
  INV_X1    g0233(.A(new_n386), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n428), .A3(new_n434), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n425), .A2(new_n429), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n382), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n253), .A2(G1), .ZN(new_n443));
  NAND2_X1  g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G270), .A3(new_n258), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n211), .A2(G45), .ZN(new_n449));
  OR2_X1    g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n444), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n266), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(G1698), .C1(new_n393), .C2(new_n394), .ZN(new_n454));
  OAI211_X1 g0254(.A(G257), .B(new_n360), .C1(new_n393), .C2(new_n394), .ZN(new_n455));
  INV_X1    g0255(.A(G303), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n278), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n282), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n211), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n304), .A2(new_n460), .A3(new_n221), .A4(new_n301), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n383), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n301), .A2(new_n221), .B1(G20), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n212), .C1(G33), .C2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT20), .B1(new_n466), .B2(new_n469), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n463), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n459), .A2(new_n473), .A3(G169), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n473), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n453), .A2(new_n458), .A3(G190), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n448), .A2(new_n452), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n282), .B2(new_n457), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n478), .C1(new_n480), .C2(new_n426), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n459), .A2(new_n473), .A3(KEYINPUT21), .A4(G169), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(G179), .A3(new_n473), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  OAI21_X1  g0286(.A(G250), .B1(new_n253), .B2(G1), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT80), .B1(new_n282), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n258), .A2(new_n489), .A3(G250), .A4(new_n449), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n488), .A2(new_n490), .B1(G274), .B2(new_n443), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(G1698), .C1(new_n393), .C2(new_n394), .ZN(new_n492));
  OAI211_X1 g0292(.A(G238), .B(new_n360), .C1(new_n393), .C2(new_n394), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n282), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n486), .B1(new_n497), .B2(G179), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n491), .A2(new_n496), .A3(KEYINPUT81), .A4(new_n251), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n290), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n372), .A2(new_n383), .ZN(new_n501));
  AOI21_X1  g0301(.A(G20), .B1(new_n273), .B2(new_n274), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G68), .ZN(new_n503));
  NAND3_X1  g0303(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n212), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n209), .B2(G87), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n297), .B2(new_n468), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n501), .B1(new_n509), .B2(new_n302), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n461), .A2(new_n372), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n491), .A2(new_n496), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n461), .A2(new_n516), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n501), .B(new_n517), .C1(new_n509), .C2(new_n302), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n497), .A2(G200), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G250), .B(new_n360), .C1(new_n393), .C2(new_n394), .ZN(new_n522));
  OAI211_X1 g0322(.A(G257), .B(G1698), .C1(new_n393), .C2(new_n394), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n282), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n447), .A2(G264), .A3(new_n258), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n452), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n528), .A2(G179), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n290), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n494), .A2(G20), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT82), .B1(new_n212), .B2(G107), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT23), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT82), .B(new_n534), .C1(new_n212), .C2(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n502), .B2(G87), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n212), .B(G87), .C1(new_n393), .C2(new_n394), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT24), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n502), .A2(new_n537), .A3(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT24), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n536), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n387), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n304), .B2(G107), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n304), .A2(new_n549), .A3(G107), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n551), .A2(new_n552), .B1(new_n362), .B2(new_n461), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n529), .B(new_n530), .C1(new_n548), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n528), .A2(new_n426), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n526), .A2(new_n527), .A3(new_n355), .A4(new_n452), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n545), .A2(new_n546), .A3(new_n536), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n546), .B1(new_n545), .B2(new_n536), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n302), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n553), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n485), .A2(new_n521), .A3(new_n554), .A4(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n275), .A2(G244), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n467), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n275), .B2(G244), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n282), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n447), .A2(new_n258), .ZN(new_n571));
  INV_X1    g0371(.A(G257), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n452), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n355), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n278), .A2(G244), .A3(new_n360), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n564), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(new_n566), .A3(new_n567), .A4(new_n467), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n573), .B1(new_n578), .B2(new_n282), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(G200), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n304), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n462), .B2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n412), .A2(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  AND2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(new_n208), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n362), .A2(KEYINPUT6), .A3(G97), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n212), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n296), .A2(new_n277), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT77), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT77), .ZN(new_n591));
  INV_X1    g0391(.A(new_n589), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n212), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n583), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT78), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(new_n302), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n595), .B2(new_n302), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n580), .B(new_n582), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n582), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n302), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT78), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n596), .A3(new_n302), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n570), .A2(new_n574), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n290), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n579), .A2(new_n251), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n599), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n563), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n442), .A2(new_n610), .ZN(G372));
  AND2_X1   g0411(.A1(new_n425), .A2(new_n437), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n353), .A2(new_n376), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n356), .A2(new_n429), .A3(new_n440), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n321), .A2(new_n323), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n310), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n442), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n582), .B1(new_n597), .B2(new_n598), .ZN(new_n619));
  INV_X1    g0419(.A(new_n608), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n513), .A2(new_n520), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n510), .A2(new_n511), .B1(new_n497), .B2(new_n290), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n514), .A2(new_n251), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n520), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n619), .A2(new_n627), .A3(new_n620), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(KEYINPUT26), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n554), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n476), .A2(new_n482), .A3(new_n483), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n627), .B(new_n562), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n626), .B1(new_n632), .B2(new_n609), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n617), .B1(new_n618), .B2(new_n634), .ZN(G369));
  NAND2_X1  g0435(.A1(new_n325), .A2(new_n212), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(G213), .ZN(new_n639));
  XOR2_X1   g0439(.A(KEYINPUT83), .B(G343), .Z(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n477), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n484), .B2(new_n643), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n641), .B1(new_n548), .B2(new_n553), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n554), .A2(new_n562), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n554), .B2(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n631), .A2(new_n642), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n630), .B2(new_n642), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(G399));
  NOR2_X1   g0455(.A1(new_n215), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n220), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n642), .B1(new_n629), .B2(new_n633), .ZN(new_n664));
  XOR2_X1   g0464(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n521), .A2(new_n619), .A3(new_n668), .A4(new_n620), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT29), .B(new_n642), .C1(new_n670), .C2(new_n633), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n480), .A2(G179), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n491), .A2(new_n496), .A3(new_n526), .A4(new_n527), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n673), .A2(new_n605), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n514), .A2(new_n480), .A3(G179), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n605), .A2(new_n528), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n676), .A2(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(KEYINPUT30), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n642), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n554), .A2(new_n562), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n683), .A2(new_n484), .A3(new_n622), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n621), .A3(new_n599), .A4(new_n642), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n685), .B2(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n641), .A2(KEYINPUT31), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n679), .A2(new_n678), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n675), .B2(KEYINPUT30), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n690));
  INV_X1    g0490(.A(new_n681), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n689), .B2(KEYINPUT85), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(G330), .B1(new_n686), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n672), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n663), .B1(new_n696), .B2(G1), .ZN(G364));
  NOR2_X1   g0497(.A1(new_n215), .A2(new_n395), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n698), .A2(G355), .B1(new_n464), .B2(new_n215), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n215), .A2(new_n278), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n660), .B2(G45), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n249), .A2(new_n253), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G13), .A2(G33), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT87), .Z(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n221), .B1(G20), .B2(new_n290), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n214), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n211), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n656), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n251), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(G20), .A2(G190), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n251), .A2(new_n426), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n212), .A2(G190), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g0522(.A(KEYINPUT33), .B(G317), .ZN(new_n723));
  AOI22_X1  g0523(.A1(G322), .A2(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n426), .A2(G179), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n725), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT89), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G283), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n724), .B1(new_n456), .B2(new_n726), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n721), .A2(new_n715), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G179), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n721), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(G311), .A2(new_n733), .B1(new_n736), .B2(G329), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n716), .A2(new_n251), .A3(new_n426), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n278), .B1(G326), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n212), .B1(new_n734), .B2(G190), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n737), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT88), .B(KEYINPUT32), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  OR3_X1    g0544(.A1(new_n735), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n395), .B1(G50), .B2(new_n738), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n743), .B1(new_n735), .B2(new_n744), .ZN(new_n747));
  INV_X1    g0547(.A(new_n741), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G97), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n728), .A2(G107), .ZN(new_n751));
  INV_X1    g0551(.A(new_n726), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G87), .A2(new_n752), .B1(new_n722), .B2(G68), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n733), .A2(G77), .B1(new_n719), .B2(G58), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n731), .A2(new_n742), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n714), .B1(new_n756), .B2(new_n707), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n709), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT90), .ZN(new_n759));
  INV_X1    g0559(.A(new_n706), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n645), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n647), .A2(new_n713), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n645), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(G396));
  NAND2_X1  g0565(.A1(new_n377), .A2(new_n642), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n380), .A2(new_n378), .B1(new_n379), .B2(new_n641), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(new_n377), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n664), .A2(new_n768), .ZN(new_n769));
  MUX2_X1   g0569(.A(new_n641), .B(new_n767), .S(new_n376), .Z(new_n770));
  OAI211_X1 g0570(.A(new_n642), .B(new_n770), .C1(new_n629), .C2(new_n633), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n713), .B1(new_n772), .B2(new_n694), .ZN(new_n773));
  INV_X1    g0573(.A(new_n694), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(new_n769), .A3(new_n771), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n722), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n777), .A2(new_n730), .B1(new_n732), .B2(new_n464), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT91), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(G303), .B2(new_n738), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT92), .Z(new_n782));
  NAND2_X1  g0582(.A1(new_n728), .A2(G87), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G294), .A2(new_n719), .B1(new_n736), .B2(G311), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(new_n749), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n395), .B1(new_n726), .B2(new_n362), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT93), .Z(new_n787));
  NOR3_X1   g0587(.A1(new_n782), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n722), .A2(G150), .B1(new_n738), .B2(G137), .ZN(new_n789));
  INV_X1    g0589(.A(G143), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n790), .B2(new_n718), .C1(new_n744), .C2(new_n732), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n728), .A2(G68), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  INV_X1    g0594(.A(G50), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n278), .B1(new_n735), .B2(new_n794), .C1(new_n795), .C2(new_n726), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G58), .B2(new_n748), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n707), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n707), .A2(new_n704), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n713), .C1(G77), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n705), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n768), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n776), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G384));
  INV_X1    g0607(.A(new_n593), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT35), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT35), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n809), .A2(new_n810), .A3(G116), .A4(new_n222), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT36), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n660), .A2(new_n277), .A3(new_n389), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n795), .B2(G68), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n214), .A2(G1), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n414), .B1(new_n430), .B2(new_n431), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n416), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n386), .B1(new_n408), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n438), .B1(new_n818), .B2(new_n639), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n424), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT37), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n433), .A2(new_n434), .ZN(new_n822));
  INV_X1    g0622(.A(new_n424), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n639), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n438), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n818), .A2(new_n639), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n821), .A2(new_n828), .B1(new_n441), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT97), .B1(new_n830), .B2(KEYINPUT38), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n824), .A2(new_n826), .A3(new_n438), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n639), .B1(new_n433), .B2(new_n434), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT96), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n833), .B(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n441), .A2(new_n834), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n686), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n353), .B(new_n356), .C1(new_n336), .C2(new_n642), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n351), .A2(new_n352), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n337), .A3(new_n641), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n768), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n830), .A2(KEYINPUT97), .A3(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n840), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n821), .A2(new_n828), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n441), .A2(new_n829), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n832), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT38), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT40), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n851), .A2(KEYINPUT40), .B1(new_n849), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT31), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n610), .B2(new_n642), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n841), .B1(new_n860), .B2(new_n682), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n442), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(G330), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT39), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT97), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n856), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n433), .A2(new_n434), .A3(new_n428), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n435), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT96), .B1(new_n418), .B2(new_n639), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n826), .A2(new_n870), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n833), .A2(new_n836), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n441), .A2(new_n834), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT38), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n866), .B(new_n850), .C1(new_n868), .C2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n845), .A2(new_n337), .A3(new_n642), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT95), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n612), .A2(new_n825), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n855), .A2(new_n856), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n844), .A2(new_n846), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n771), .B2(new_n766), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n442), .A2(new_n671), .A3(new_n666), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n617), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n888), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n865), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n211), .B2(new_n710), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n865), .A2(new_n891), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n812), .B1(new_n814), .B2(new_n815), .C1(new_n893), .C2(new_n894), .ZN(G367));
  INV_X1    g0695(.A(new_n700), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n240), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n708), .B1(new_n216), .B2(new_n372), .ZN(new_n898));
  INV_X1    g0698(.A(new_n738), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n790), .B1(new_n726), .B2(new_n202), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n395), .B(new_n900), .C1(G150), .C2(new_n719), .ZN(new_n901));
  INV_X1    g0701(.A(new_n727), .ZN(new_n902));
  AOI22_X1  g0702(.A1(G77), .A2(new_n902), .B1(new_n736), .B2(G137), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n733), .A2(G50), .B1(new_n722), .B2(G159), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n748), .A2(G68), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n733), .A2(G283), .B1(new_n738), .B2(G311), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n278), .B1(new_n736), .B2(G317), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n907), .B(new_n908), .C1(new_n362), .C2(new_n741), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n752), .A2(G116), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT46), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n902), .A2(G97), .B1(new_n719), .B2(G303), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n911), .B(new_n912), .C1(new_n740), .C2(new_n777), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n906), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT47), .Z(new_n915));
  INV_X1    g0715(.A(new_n707), .ZN(new_n916));
  OAI221_X1 g0716(.A(new_n713), .B1(new_n897), .B2(new_n898), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT105), .ZN(new_n918));
  INV_X1    g0718(.A(new_n518), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n624), .A2(new_n919), .A3(new_n625), .A4(new_n641), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT98), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n627), .B1(new_n518), .B2(new_n642), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n920), .A2(new_n921), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n760), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT100), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n621), .B(new_n599), .C1(new_n604), .C2(new_n642), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n621), .B2(new_n642), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n931), .A2(new_n653), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT42), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n930), .A2(new_n554), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n934), .A2(new_n621), .ZN(new_n935));
  OAI221_X1 g0735(.A(new_n929), .B1(new_n932), .B2(new_n933), .C1(new_n935), .C2(new_n641), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n641), .B1(new_n934), .B2(new_n621), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT100), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n936), .A2(new_n939), .B1(new_n933), .B2(new_n932), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n925), .B2(KEYINPUT99), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(KEYINPUT99), .B2(new_n925), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT101), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n940), .A2(new_n949), .A3(new_n943), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(new_n940), .B2(new_n943), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n651), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n931), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n940), .A2(new_n943), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT101), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n940), .A2(new_n949), .A3(new_n943), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(new_n954), .A3(new_n948), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n956), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n931), .A2(new_n654), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n931), .A2(new_n654), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n953), .A2(KEYINPUT103), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n653), .ZN(new_n973));
  INV_X1    g0773(.A(new_n652), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n650), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n647), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n672), .A2(new_n694), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n966), .A2(new_n970), .A3(new_n968), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n972), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(new_n696), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n656), .B(KEYINPUT41), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n711), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n962), .A2(new_n963), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n963), .B1(new_n962), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n928), .B1(new_n984), .B2(new_n985), .ZN(G387));
  NOR2_X1   g0786(.A1(new_n977), .A2(new_n657), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n696), .B2(new_n976), .ZN(new_n988));
  INV_X1    g0788(.A(new_n658), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n989), .A2(new_n698), .B1(new_n362), .B2(new_n215), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n237), .A2(new_n253), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n298), .A2(new_n795), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n658), .B(new_n253), .C1(new_n203), .C2(new_n277), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n700), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n990), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n714), .B1(new_n996), .B2(new_n708), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n650), .B2(new_n760), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n722), .A2(G311), .B1(new_n738), .B2(G322), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n732), .A2(new_n456), .B1(new_n718), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT107), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT108), .Z(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G294), .A2(new_n752), .B1(new_n748), .B2(G283), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n727), .A2(new_n464), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n278), .B(new_n1013), .C1(G326), .C2(new_n736), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n726), .A2(new_n277), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n395), .B(new_n1016), .C1(G150), .C2(new_n736), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n468), .B2(new_n729), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT106), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n777), .A2(new_n299), .B1(new_n795), .B2(new_n718), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n899), .A2(new_n744), .B1(new_n732), .B2(new_n203), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n741), .A2(new_n372), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1015), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n998), .B1(new_n1024), .B2(new_n707), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n712), .B2(new_n976), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n988), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT109), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(G393));
  XNOR2_X1  g0830(.A(new_n969), .B(new_n651), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n656), .B(new_n979), .C1(new_n1031), .C2(new_n977), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n712), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n395), .B1(new_n752), .B2(G68), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n783), .B(new_n1034), .C1(new_n790), .C2(new_n735), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n719), .A2(G159), .B1(new_n738), .B2(G150), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT51), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n748), .A2(G77), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n299), .B2(new_n732), .C1(new_n777), .C2(new_n795), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n719), .A2(G311), .B1(new_n738), .B2(G317), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n751), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n736), .A2(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n740), .B2(new_n732), .C1(new_n777), .C2(new_n456), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n395), .B1(new_n741), .B2(new_n464), .C1(new_n730), .C2(new_n726), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n707), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n708), .B1(new_n468), .B2(new_n216), .C1(new_n245), .C2(new_n896), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT110), .Z(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n1052), .A3(new_n713), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT112), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n760), .B2(new_n931), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1032), .A2(new_n1033), .A3(new_n1055), .ZN(G390));
  NAND2_X1  g0856(.A1(new_n774), .A2(new_n847), .ZN(new_n1057));
  AND4_X1   g0857(.A1(KEYINPUT97), .A2(new_n852), .A3(new_n853), .A4(KEYINPUT38), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n831), .B2(new_n839), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n767), .A2(new_n377), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n642), .B(new_n1060), .C1(new_n670), .C2(new_n633), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n766), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n879), .B1(new_n1062), .B2(new_n884), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1059), .B2(new_n866), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n886), .A2(new_n879), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1057), .B(new_n1064), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n847), .B(G330), .C1(new_n686), .C2(new_n842), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT113), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT113), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n861), .A2(new_n1071), .A3(G330), .A4(new_n847), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n879), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n771), .A2(new_n766), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n884), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n877), .A2(new_n880), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1068), .A2(new_n1079), .A3(new_n712), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n861), .A2(G330), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n889), .B(new_n617), .C1(new_n618), .C2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(G330), .B(new_n770), .C1(new_n686), .C2(new_n693), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n885), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1070), .A2(new_n1087), .A3(new_n1072), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1062), .B1(new_n774), .B2(new_n847), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n885), .B1(new_n1084), .B2(new_n768), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1088), .A2(new_n1075), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1083), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1075), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1085), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n1068), .A3(new_n1079), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n656), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n278), .B1(new_n727), .B2(new_n795), .ZN(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1098), .A2(KEYINPUT115), .B1(new_n1099), .B2(new_n735), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT115), .B2(new_n1098), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT116), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G132), .A2(new_n719), .B1(new_n722), .B2(G137), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n733), .A2(new_n1105), .B1(new_n738), .B2(G128), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n752), .A2(G150), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G159), .B2(new_n748), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1102), .A2(new_n1103), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n777), .A2(new_n362), .B1(new_n735), .B2(new_n740), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n278), .B(new_n1111), .C1(G87), .C2(new_n752), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n899), .A2(new_n730), .B1(new_n718), .B2(new_n464), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G97), .B2(new_n733), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1112), .A2(new_n793), .A3(new_n1039), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n916), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n714), .B(new_n1116), .C1(new_n299), .C2(new_n800), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1066), .B2(new_n705), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1082), .A2(new_n1097), .A3(new_n1118), .ZN(G378));
  NAND2_X1  g0919(.A1(new_n308), .A2(new_n825), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n324), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n324), .A2(new_n1120), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n881), .A2(new_n887), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n881), .B2(new_n887), .ZN(new_n1129));
  INV_X1    g0929(.A(G330), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n858), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n888), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n851), .A2(KEYINPUT40), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT40), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n849), .A2(new_n1135), .A3(new_n883), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1130), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n881), .A2(new_n887), .A3(new_n1127), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1085), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1096), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n657), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT57), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT118), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1140), .A2(new_n1142), .A3(new_n1148), .A4(KEYINPUT57), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1132), .A2(new_n803), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n713), .B1(G50), .B2(new_n801), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n777), .A2(new_n794), .B1(new_n1099), .B2(new_n899), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G137), .A2(new_n733), .B1(new_n752), .B2(new_n1105), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n718), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1153), .B(new_n1156), .C1(G150), .C2(new_n748), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n736), .C2(G124), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n744), .B2(new_n727), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT117), .Z(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n727), .A2(new_n202), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G283), .B2(new_n736), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1016), .A2(G41), .A3(new_n278), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n905), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n899), .A2(new_n464), .B1(new_n732), .B2(new_n372), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n777), .A2(new_n468), .B1(new_n362), .B2(new_n718), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n795), .B1(new_n393), .B2(G41), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1164), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1152), .B1(new_n1175), .B2(new_n707), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1140), .A2(new_n712), .B1(new_n1151), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1150), .A2(new_n1177), .ZN(G375));
  OAI22_X1  g0978(.A1(new_n726), .A2(new_n744), .B1(new_n735), .B2(new_n1155), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT121), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n395), .B(new_n1165), .C1(G50), .C2(new_n748), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n719), .A2(G137), .B1(new_n738), .B2(G132), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G150), .A2(new_n733), .B1(new_n722), .B2(new_n1105), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n777), .A2(new_n464), .B1(new_n732), .B2(new_n362), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n278), .B(new_n1185), .C1(G294), .C2(new_n738), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n726), .A2(new_n468), .B1(new_n735), .B2(new_n456), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT119), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(new_n277), .C2(new_n729), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1022), .B1(G283), .B2(new_n719), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT120), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1184), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n707), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n713), .C1(G68), .C2(new_n801), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n885), .B2(new_n704), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1091), .B2(new_n711), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1095), .A2(new_n981), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1091), .A2(new_n1085), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1199), .B2(new_n1201), .ZN(G381));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1150), .A2(new_n1203), .A3(new_n1177), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1028), .A2(new_n764), .A3(new_n1029), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1205), .A2(G384), .A3(G390), .ZN(new_n1206));
  OR4_X1    g1006(.A1(G387), .A2(new_n1204), .A3(new_n1206), .A4(G381), .ZN(G407));
  NAND2_X1  g1007(.A1(new_n640), .A2(G213), .ZN(new_n1208));
  OAI211_X1 g1008(.A(G407), .B(G213), .C1(new_n1204), .C2(new_n1208), .ZN(G409));
  INV_X1    g1009(.A(KEYINPUT124), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1205), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1210), .A3(new_n1205), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n954), .B1(new_n960), .B2(new_n948), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n955), .B(new_n947), .C1(new_n958), .C2(new_n959), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n982), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT104), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n983), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G390), .B1(new_n1220), .B2(new_n928), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n927), .B(new_n1222), .C1(new_n1219), .C2(new_n983), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1215), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G387), .A2(new_n1222), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1214), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(new_n1212), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1220), .A2(new_n928), .A3(G390), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1224), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G375), .A2(G378), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1143), .A2(new_n981), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1177), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1208), .C1(G378), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT60), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1200), .B1(new_n1095), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1091), .A2(KEYINPUT60), .A3(new_n1085), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n656), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(KEYINPUT122), .A3(new_n656), .A4(new_n1237), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1197), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(G384), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1234), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1230), .B1(KEYINPUT63), .B2(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1244), .A2(KEYINPUT63), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1242), .B(new_n806), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n640), .A2(G213), .A3(G2897), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT123), .Z(new_n1250));
  OR2_X1    g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1234), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1247), .B(new_n1253), .C1(new_n1244), .C2(new_n1255), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1234), .A2(KEYINPUT62), .A3(new_n1243), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1230), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1254), .A2(new_n1258), .ZN(G405));
  AND3_X1   g1059(.A1(new_n1150), .A2(new_n1203), .A3(new_n1177), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1203), .B1(new_n1150), .B2(new_n1177), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1243), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1243), .B(KEYINPUT126), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1231), .A2(new_n1204), .A3(new_n1248), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT125), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1231), .A2(new_n1248), .A3(new_n1269), .A4(new_n1204), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1271), .A3(new_n1230), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1266), .A2(new_n1271), .A3(new_n1230), .A4(KEYINPUT127), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1230), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1278), .ZN(G402));
endmodule


