//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n444, new_n445, new_n446, new_n448, new_n452,
    new_n453, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g024(.A(G452), .Z(G391));
  AND2_X1   g025(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g029(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g030(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g031(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT2), .Z(new_n458));
  NAND4_X1  g033(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(new_n461), .ZN(G261));
  INV_X1    g037(.A(G261), .ZN(G325));
  NAND2_X1  g038(.A1(new_n460), .A2(G567), .ZN(new_n464));
  INV_X1    g039(.A(G2106), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT70), .B1(new_n468), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT71), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n469), .A2(new_n472), .A3(new_n476), .A4(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n480), .A2(new_n482), .A3(G137), .A4(new_n471), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G137), .A4(new_n471), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n478), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G160));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n483), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n489), .A2(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G124), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n496), .A2(new_n497), .A3(new_n471), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G136), .ZN(new_n503));
  OR2_X1    g078(.A1(G100), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n500), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G162));
  NAND4_X1  g082(.A1(new_n480), .A2(new_n482), .A3(G138), .A4(new_n471), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G114), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n513), .A2(new_n468), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n489), .B2(G126), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n515), .B2(new_n471), .ZN(new_n516));
  INV_X1    g091(.A(G138), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n489), .A2(new_n510), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G102), .A2(G2104), .ZN(new_n520));
  AOI21_X1  g095(.A(G2105), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G164));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n529), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n525), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n536), .B(new_n540), .C1(new_n525), .C2(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT5), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n544), .A2(new_n546), .A3(G63), .A4(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n523), .A2(KEYINPUT74), .A3(G63), .A4(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g126(.A1(KEYINPUT6), .A2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(KEYINPUT6), .A2(G651), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G51), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n551), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT75), .B1(new_n551), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n542), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n542), .B(KEYINPUT77), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(G168));
  INV_X1    g137(.A(G90), .ZN(new_n563));
  INV_X1    g138(.A(G52), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n525), .A2(new_n563), .B1(new_n527), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT78), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n565), .B1(new_n567), .B2(G651), .ZN(G171));
  INV_X1    g143(.A(G81), .ZN(new_n569));
  INV_X1    g144(.A(G43), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n525), .A2(new_n569), .B1(new_n527), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n531), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G188));
  NAND3_X1  g155(.A1(new_n524), .A2(KEYINPUT79), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT9), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n554), .A2(KEYINPUT79), .A3(new_n584), .A4(G53), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n531), .ZN(new_n588));
  INV_X1    g163(.A(new_n525), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G91), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n583), .A2(new_n585), .B1(G91), .B2(new_n589), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n588), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G299));
  INV_X1    g171(.A(G171), .ZN(G301));
  INV_X1    g172(.A(G168), .ZN(G286));
  NAND3_X1  g173(.A1(new_n589), .A2(KEYINPUT81), .A3(G87), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  INV_X1    g175(.A(G87), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n525), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  INV_X1    g179(.A(G49), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n527), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n554), .A2(KEYINPUT82), .A3(G49), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n523), .A2(G74), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n606), .A2(new_n607), .B1(G651), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n603), .A2(new_n609), .ZN(G288));
  INV_X1    g185(.A(G86), .ZN(new_n611));
  INV_X1    g186(.A(G48), .ZN(new_n612));
  OAI22_X1  g187(.A1(new_n525), .A2(new_n611), .B1(new_n527), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n531), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(G305));
  INV_X1    g192(.A(G85), .ZN(new_n618));
  INV_X1    g193(.A(G47), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n525), .A2(new_n618), .B1(new_n527), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(new_n531), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n620), .A2(new_n622), .ZN(G290));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT83), .B1(new_n525), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n523), .A2(new_n524), .A3(new_n626), .A4(G92), .ZN(new_n627));
  AOI21_X1  g202(.A(KEYINPUT10), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n523), .A2(G66), .ZN(new_n630));
  INV_X1    g205(.A(G79), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n543), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n632), .A2(G651), .B1(G54), .B2(new_n554), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(G171), .ZN(G321));
  XOR2_X1   g213(.A(G321), .B(KEYINPUT84), .Z(G284));
  NAND2_X1  g214(.A1(G299), .A2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G297));
  OAI21_X1  g216(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G280));
  INV_X1    g217(.A(new_n635), .ZN(new_n643));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(G860), .ZN(G148));
  OAI21_X1  g220(.A(KEYINPUT85), .B1(new_n574), .B2(G868), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G868), .ZN(new_n648));
  MUX2_X1   g223(.A(KEYINPUT85), .B(new_n646), .S(new_n648), .Z(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g225(.A(new_n473), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n489), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n499), .A2(G123), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n502), .A2(G135), .ZN(new_n657));
  OR2_X1    g232(.A1(G99), .A2(G2105), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n658), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2435), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2438), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT14), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1341), .B(G1348), .Z(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n673), .B(new_n676), .Z(new_n677));
  AND2_X1   g252(.A1(new_n677), .A2(G14), .ZN(G401));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT90), .Z(new_n681));
  XNOR2_X1  g256(.A(G2072), .B(G2078), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT91), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(KEYINPUT92), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT17), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n686), .C1(new_n681), .C2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n681), .A2(new_n685), .A3(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n680), .A2(new_n685), .A3(new_n682), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT18), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2096), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2100), .Z(G227));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n697), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n699), .A2(new_n701), .A3(new_n703), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n706), .B(new_n707), .C1(new_n705), .C2(new_n704), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(G1986), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(G229));
  NOR2_X1   g289(.A1(G16), .A2(G22), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G166), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT95), .B(G1971), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT94), .B1(G16), .B2(G23), .ZN(new_n719));
  OR3_X1    g294(.A1(KEYINPUT94), .A2(G16), .A3(G23), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n719), .B(new_n720), .C1(G288), .C2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(G6), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n616), .B2(new_n721), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n718), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n718), .A2(new_n724), .A3(KEYINPUT34), .A4(new_n728), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n499), .A2(G119), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n502), .A2(G131), .ZN(new_n735));
  NOR2_X1   g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT35), .B(G1991), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G24), .B(G290), .S(G16), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1986), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n733), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n733), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G35), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT103), .B1(new_n752), .B2(G29), .ZN(new_n753));
  OR3_X1    g328(.A1(new_n752), .A2(KEYINPUT103), .A3(G29), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(G162), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G2090), .ZN(new_n758));
  NAND2_X1  g333(.A1(G299), .A2(G16), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n721), .A2(KEYINPUT23), .A3(G20), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G20), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G16), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT104), .B(G1956), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(G29), .A2(G32), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n502), .A2(G141), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n499), .A2(G129), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n651), .A2(G105), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  NAND4_X1  g347(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n755), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n721), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n721), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1961), .Z(new_n779));
  NAND4_X1  g354(.A1(new_n758), .A2(new_n766), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n774), .A2(new_n775), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n782));
  INV_X1    g357(.A(new_n660), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n755), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n660), .A2(KEYINPUT100), .A3(G29), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G28), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n788), .A2(new_n789), .A3(new_n755), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n493), .A2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  INV_X1    g367(.A(G34), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(KEYINPUT24), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(KEYINPUT24), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n755), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n800));
  INV_X1    g375(.A(G139), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n799), .B1(new_n471), .B2(new_n800), .C1(new_n501), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G33), .B(new_n802), .S(G29), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(new_n444), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n786), .A2(new_n790), .A3(new_n797), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n780), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n792), .B1(new_n791), .B2(new_n796), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT98), .B(KEYINPUT28), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n755), .A2(G26), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n812));
  INV_X1    g387(.A(G128), .ZN(new_n813));
  INV_X1    g388(.A(G140), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n498), .B2(new_n813), .C1(new_n814), .C2(new_n501), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(G29), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n815), .B2(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n810), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G2067), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n807), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G4), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n643), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT96), .B(G1348), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n764), .A2(new_n765), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n757), .A2(G2090), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(G286), .A2(G16), .ZN(new_n832));
  INV_X1    g407(.A(G1966), .ZN(new_n833));
  INV_X1    g408(.A(G21), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n832), .B(new_n833), .C1(G16), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT31), .B(G11), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n806), .A2(new_n831), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n832), .B1(G16), .B2(new_n834), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G1966), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT99), .Z(new_n841));
  NOR3_X1   g416(.A1(new_n751), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n721), .A2(G19), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n574), .B2(new_n721), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1341), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G27), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT102), .B1(new_n847), .B2(G29), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n847), .A2(KEYINPUT102), .A3(G29), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(G164), .C2(new_n755), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n445), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n842), .A2(KEYINPUT105), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  INV_X1    g428(.A(new_n838), .ZN(new_n854));
  INV_X1    g429(.A(new_n841), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n854), .A2(new_n750), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n856), .B2(new_n845), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n857), .ZN(G311));
  NAND3_X1  g433(.A1(new_n842), .A2(new_n846), .A3(new_n851), .ZN(G150));
  NAND2_X1  g434(.A1(new_n554), .A2(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  OAI221_X1 g437(.A(new_n860), .B1(new_n525), .B2(new_n861), .C1(new_n862), .C2(new_n531), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  XOR2_X1   g440(.A(new_n574), .B(new_n863), .Z(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n635), .A2(new_n644), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n870), .B2(G860), .ZN(G145));
  NAND2_X1  g446(.A1(new_n499), .A2(G130), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n502), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n738), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT107), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n653), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n802), .A2(KEYINPUT106), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n802), .B(KEYINPUT106), .ZN(new_n881));
  INV_X1    g456(.A(G164), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n815), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n773), .ZN(new_n884));
  MUX2_X1   g459(.A(new_n880), .B(new_n881), .S(new_n884), .Z(new_n885));
  OR2_X1    g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n879), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n506), .B(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n660), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n890), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT40), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n892), .A2(new_n897), .A3(new_n893), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G395));
  NOR2_X1   g474(.A1(new_n863), .A2(G868), .ZN(new_n900));
  INV_X1    g475(.A(new_n866), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n647), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n594), .A2(KEYINPUT80), .A3(new_n588), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT80), .B1(new_n594), .B2(new_n588), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n635), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n634), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n628), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n593), .A2(new_n907), .A3(new_n595), .A4(new_n633), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT41), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT41), .B1(new_n905), .B2(new_n908), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n918));
  XOR2_X1   g493(.A(G303), .B(new_n918), .Z(new_n919));
  INV_X1    g494(.A(G288), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G303), .B(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G288), .ZN(new_n923));
  XNOR2_X1  g498(.A(G305), .B(G290), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n921), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n916), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n917), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n900), .B1(new_n930), .B2(G868), .ZN(G295));
  AOI21_X1  g506(.A(new_n900), .B1(new_n930), .B2(G868), .ZN(G331));
  INV_X1    g507(.A(new_n909), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n560), .A2(new_n561), .A3(G301), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G301), .B1(new_n560), .B2(new_n561), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n936), .A3(new_n901), .ZN(new_n937));
  NAND2_X1  g512(.A1(G168), .A2(G171), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n866), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n933), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n866), .A3(new_n934), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n901), .B1(new_n935), .B2(new_n936), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n913), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n943), .A3(new_n927), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n943), .A3(new_n927), .A4(KEYINPUT112), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n927), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n913), .A2(new_n941), .A3(new_n942), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n909), .B1(new_n942), .B2(new_n941), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT111), .A3(new_n893), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n927), .B1(new_n940), .B2(new_n943), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(G37), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n948), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n948), .A2(new_n958), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n516), .B2(new_n521), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n478), .A2(G40), .A3(new_n486), .A4(new_n492), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n738), .B(new_n741), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT115), .Z(new_n976));
  XOR2_X1   g551(.A(new_n773), .B(G1996), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n815), .B(new_n820), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n974), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n981), .A2(new_n973), .A3(new_n972), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT48), .Z(new_n983));
  OR2_X1    g558(.A1(new_n738), .A2(new_n741), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n979), .A2(new_n984), .B1(G2067), .B2(new_n815), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n980), .A2(new_n983), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n978), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n974), .B1(new_n987), .B2(new_n773), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n972), .A2(G1996), .A3(new_n973), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(KEYINPUT46), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(KEYINPUT46), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n986), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n973), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n969), .C1(new_n516), .C2(new_n521), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n972), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n972), .A2(new_n996), .A3(KEYINPUT116), .A4(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT117), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(G1971), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n970), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT50), .B(new_n969), .C1(new_n516), .C2(new_n521), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n996), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(G2090), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(new_n1008), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G166), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT55), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT118), .B(KEYINPUT119), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(KEYINPUT55), .A3(new_n1019), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(new_n1022), .C1(KEYINPUT55), .C2(new_n1017), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1015), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  OAI221_X1 g600(.A(G8), .B1(new_n973), .B2(new_n970), .C1(G288), .C2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(G1976), .B2(new_n920), .ZN(new_n1028));
  OR2_X1    g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G305), .A2(G1981), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n970), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1016), .B1(new_n1034), .B2(new_n996), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1026), .A2(KEYINPUT120), .A3(KEYINPUT52), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT120), .B1(new_n1026), .B2(KEYINPUT52), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1028), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1024), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n973), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n792), .A2(new_n1043), .B1(new_n998), .B2(new_n833), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(G286), .A3(new_n1016), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1016), .B1(new_n1046), .B2(new_n1014), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1047), .B2(new_n1023), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT63), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1041), .A2(new_n1015), .A3(G8), .A4(new_n1023), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1037), .A2(new_n1025), .A3(new_n920), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1029), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1035), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT121), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1050), .A2(KEYINPUT121), .A3(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1044), .A2(new_n1016), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G286), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT125), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1044), .A2(G168), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT126), .A2(KEYINPUT51), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1000), .A2(new_n445), .A3(new_n1001), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(G2078), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n972), .A2(new_n996), .A3(new_n997), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1043), .B2(G1961), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G301), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1076), .A2(KEYINPUT62), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1068), .A2(new_n1077), .B1(new_n1078), .B2(new_n1045), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n972), .A2(new_n996), .A3(new_n997), .A4(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT122), .B(G1956), .Z(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1043), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n591), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n594), .A2(KEYINPUT57), .A3(new_n588), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1034), .A2(new_n996), .A3(new_n820), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1043), .B2(G1348), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n643), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1090), .B(new_n1084), .C1(new_n1043), .C2(new_n1085), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1085), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1013), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1090), .B1(new_n1104), .B2(new_n1084), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1098), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1102), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT124), .B(new_n1102), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n635), .B(new_n1093), .C1(new_n1043), .C2(G1348), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1095), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n970), .B2(new_n973), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n998), .B2(G1996), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n574), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1120), .A3(new_n574), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n635), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1114), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1101), .B1(new_n1111), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1071), .A2(G301), .A3(new_n1075), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1081), .A2(KEYINPUT54), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n1129));
  AOI211_X1 g704(.A(G171), .B(new_n1074), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1076), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1082), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1079), .B1(new_n1133), .B2(new_n1068), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1014), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1023), .B1(new_n1136), .B2(G8), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1042), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1056), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n981), .A2(KEYINPUT113), .A3(new_n1140), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n974), .C1(KEYINPUT113), .C2(new_n1140), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT114), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n980), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n995), .B1(new_n1139), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g720(.A(G319), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G229), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g722(.A1(G401), .A2(G227), .ZN(new_n1149));
  AND4_X1   g723(.A1(new_n895), .A2(new_n965), .A3(new_n1148), .A4(new_n1149), .ZN(G308));
  NAND4_X1  g724(.A1(new_n895), .A2(new_n965), .A3(new_n1148), .A4(new_n1149), .ZN(G225));
endmodule


