

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758;

  INV_X1 U364 ( .A(n660), .ZN(n342) );
  INV_X1 U365 ( .A(KEYINPUT56), .ZN(n344) );
  AND2_X1 U366 ( .A1(n376), .A2(n377), .ZN(n375) );
  XNOR2_X1 U367 ( .A(n612), .B(n611), .ZN(n620) );
  NOR2_X1 U368 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U369 ( .A(n542), .B(n541), .ZN(n610) );
  NAND2_X1 U370 ( .A1(n538), .A2(n349), .ZN(n542) );
  OR2_X1 U371 ( .A1(n371), .A2(n370), .ZN(n519) );
  XNOR2_X1 U372 ( .A(n393), .B(n511), .ZN(n515) );
  XNOR2_X1 U373 ( .A(n473), .B(n413), .ZN(n586) );
  XNOR2_X1 U374 ( .A(n501), .B(G134), .ZN(n473) );
  XNOR2_X1 U375 ( .A(n415), .B(n414), .ZN(n495) );
  XNOR2_X1 U376 ( .A(G116), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U377 ( .A(n343), .B(n342), .ZN(G57) );
  NAND2_X1 U378 ( .A1(n659), .A2(n668), .ZN(n343) );
  XNOR2_X1 U379 ( .A(n345), .B(n344), .ZN(G51) );
  NAND2_X1 U380 ( .A1(n669), .A2(n668), .ZN(n345) );
  XNOR2_X1 U381 ( .A(n596), .B(n595), .ZN(n379) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n483) );
  INV_X1 U383 ( .A(n608), .ZN(n599) );
  INV_X2 U384 ( .A(G953), .ZN(n454) );
  XNOR2_X2 U385 ( .A(n467), .B(KEYINPUT79), .ZN(n557) );
  XNOR2_X2 U386 ( .A(n562), .B(KEYINPUT41), .ZN(n719) );
  NOR2_X1 U387 ( .A1(n525), .A2(n450), .ZN(n391) );
  INV_X1 U388 ( .A(KEYINPUT64), .ZN(n398) );
  XNOR2_X1 U389 ( .A(n399), .B(n398), .ZN(n397) );
  NAND2_X1 U390 ( .A1(n388), .A2(n350), .ZN(n399) );
  AND2_X1 U391 ( .A1(n407), .A2(n635), .ZN(n410) );
  NOR2_X1 U392 ( .A1(n619), .A2(n618), .ZN(n631) );
  NAND2_X1 U393 ( .A1(n400), .A2(n583), .ZN(n634) );
  XNOR2_X1 U394 ( .A(n601), .B(n600), .ZN(n718) );
  XNOR2_X1 U395 ( .A(n391), .B(n390), .ZN(n546) );
  XNOR2_X1 U396 ( .A(n392), .B(n446), .ZN(n525) );
  XNOR2_X1 U397 ( .A(n476), .B(n671), .ZN(n554) );
  OR2_X1 U398 ( .A1(n656), .A2(G902), .ZN(n422) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT15), .ZN(n633) );
  XNOR2_X1 U400 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n433) );
  XNOR2_X1 U401 ( .A(G128), .B(G119), .ZN(n435) );
  OR2_X1 U402 ( .A1(G953), .A2(G952), .ZN(n427) );
  NOR2_X1 U403 ( .A1(n564), .A2(n528), .ZN(n568) );
  XNOR2_X1 U404 ( .A(KEYINPUT90), .B(KEYINPUT0), .ZN(n520) );
  NAND2_X1 U405 ( .A1(n519), .A2(n518), .ZN(n521) );
  NAND2_X1 U406 ( .A1(n379), .A2(n378), .ZN(n374) );
  AND2_X1 U407 ( .A1(n346), .A2(KEYINPUT88), .ZN(n378) );
  NAND2_X1 U408 ( .A1(n514), .A2(n348), .ZN(n372) );
  NAND2_X1 U409 ( .A1(n597), .A2(n527), .ZN(n564) );
  OR2_X2 U410 ( .A1(n637), .A2(G902), .ZN(n392) );
  XNOR2_X1 U411 ( .A(n565), .B(n530), .ZN(n385) );
  XNOR2_X1 U412 ( .A(n358), .B(n401), .ZN(n400) );
  XNOR2_X1 U413 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  NAND2_X1 U414 ( .A1(n631), .A2(n630), .ZN(n389) );
  XNOR2_X1 U415 ( .A(n586), .B(G146), .ZN(n459) );
  NAND2_X1 U416 ( .A1(n507), .A2(n633), .ZN(n393) );
  XNOR2_X1 U417 ( .A(n568), .B(n368), .ZN(n367) );
  INV_X1 U418 ( .A(KEYINPUT107), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n540), .B(n539), .ZN(n541) );
  BUF_X1 U420 ( .A(n385), .Z(n382) );
  AND2_X2 U421 ( .A1(n397), .A2(n356), .ZN(n641) );
  NAND2_X1 U422 ( .A1(KEYINPUT88), .A2(KEYINPUT44), .ZN(n377) );
  NAND2_X1 U423 ( .A1(n578), .A2(n577), .ZN(n357) );
  INV_X1 U424 ( .A(KEYINPUT46), .ZN(n402) );
  INV_X1 U425 ( .A(KEYINPUT2), .ZN(n409) );
  INV_X1 U426 ( .A(G237), .ZN(n423) );
  XNOR2_X1 U427 ( .A(G113), .B(KEYINPUT74), .ZN(n414) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n480) );
  XNOR2_X1 U429 ( .A(G131), .B(G140), .ZN(n479) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n477) );
  XOR2_X1 U431 ( .A(G122), .B(G104), .Z(n478) );
  NAND2_X1 U432 ( .A1(n634), .A2(n409), .ZN(n387) );
  INV_X1 U433 ( .A(n633), .ZN(n408) );
  NAND2_X1 U434 ( .A1(n636), .A2(n409), .ZN(n388) );
  NOR2_X1 U435 ( .A1(n515), .A2(n352), .ZN(n370) );
  NAND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U437 ( .A1(n563), .A2(n703), .ZN(n425) );
  XNOR2_X1 U438 ( .A(n432), .B(n386), .ZN(n470) );
  XNOR2_X1 U439 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n432) );
  XNOR2_X1 U440 ( .A(n469), .B(n468), .ZN(n472) );
  INV_X1 U441 ( .A(KEYINPUT7), .ZN(n468) );
  XNOR2_X1 U442 ( .A(n369), .B(KEYINPUT9), .ZN(n469) );
  XNOR2_X1 U443 ( .A(G107), .B(G122), .ZN(n369) );
  XNOR2_X1 U444 ( .A(G107), .B(G104), .ZN(n451) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n426) );
  NAND2_X1 U446 ( .A1(n381), .A2(n380), .ZN(n604) );
  INV_X1 U447 ( .A(n602), .ZN(n380) );
  NAND2_X1 U448 ( .A1(n384), .A2(n383), .ZN(n547) );
  INV_X1 U449 ( .A(n385), .ZN(n383) );
  NAND2_X1 U450 ( .A1(n553), .A2(n554), .ZN(n572) );
  XNOR2_X1 U451 ( .A(n405), .B(KEYINPUT28), .ZN(n404) );
  NOR2_X1 U452 ( .A1(n564), .A2(n688), .ZN(n405) );
  INV_X1 U453 ( .A(KEYINPUT100), .ZN(n595) );
  OR2_X1 U454 ( .A1(n645), .A2(G902), .ZN(n461) );
  INV_X1 U455 ( .A(KEYINPUT69), .ZN(n390) );
  BUF_X1 U456 ( .A(n563), .Z(n691) );
  BUF_X1 U457 ( .A(n536), .Z(n602) );
  NAND2_X1 U458 ( .A1(n407), .A2(n394), .ZN(n356) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n394) );
  INV_X1 U460 ( .A(KEYINPUT86), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n366), .B(KEYINPUT36), .ZN(n569) );
  NAND2_X1 U462 ( .A1(n367), .A2(n351), .ZN(n366) );
  XNOR2_X1 U463 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n611) );
  XNOR2_X1 U464 ( .A(n572), .B(n365), .ZN(n738) );
  INV_X1 U465 ( .A(KEYINPUT102), .ZN(n365) );
  NOR2_X1 U466 ( .A1(n691), .A2(n598), .ZN(n346) );
  AND2_X1 U467 ( .A1(n356), .A2(G475), .ZN(n347) );
  XOR2_X1 U468 ( .A(KEYINPUT67), .B(KEYINPUT19), .Z(n348) );
  AND2_X1 U469 ( .A1(n702), .A2(n680), .ZN(n349) );
  AND2_X1 U470 ( .A1(n387), .A2(n408), .ZN(n350) );
  NOR2_X1 U471 ( .A1(n556), .A2(n514), .ZN(n351) );
  OR2_X1 U472 ( .A1(n514), .A2(n348), .ZN(n352) );
  NOR2_X1 U473 ( .A1(n681), .A2(n382), .ZN(n353) );
  XOR2_X1 U474 ( .A(n656), .B(n657), .Z(n354) );
  XOR2_X1 U475 ( .A(n666), .B(n665), .Z(n355) );
  NAND2_X1 U476 ( .A1(n679), .A2(n356), .ZN(n725) );
  NAND2_X1 U477 ( .A1(n357), .A2(n403), .ZN(n363) );
  NAND2_X1 U478 ( .A1(n360), .A2(n359), .ZN(n358) );
  XNOR2_X1 U479 ( .A(n364), .B(n402), .ZN(n359) );
  NAND2_X1 U480 ( .A1(n363), .A2(n361), .ZN(n360) );
  NAND2_X1 U481 ( .A1(n578), .A2(n362), .ZN(n361) );
  AND2_X1 U482 ( .A1(n577), .A2(KEYINPUT72), .ZN(n362) );
  NAND2_X1 U483 ( .A1(n662), .A2(n593), .ZN(n364) );
  INV_X1 U484 ( .A(n537), .ZN(n553) );
  INV_X1 U485 ( .A(n738), .ZN(n551) );
  NAND2_X1 U486 ( .A1(n515), .A2(n348), .ZN(n373) );
  NAND2_X1 U487 ( .A1(n375), .A2(n374), .ZN(n613) );
  NAND2_X1 U488 ( .A1(n620), .A2(KEYINPUT88), .ZN(n376) );
  NAND2_X1 U489 ( .A1(n379), .A2(n346), .ZN(n622) );
  INV_X1 U490 ( .A(n718), .ZN(n381) );
  INV_X1 U491 ( .A(n683), .ZN(n384) );
  NAND2_X1 U492 ( .A1(n683), .A2(n382), .ZN(n685) );
  NAND2_X1 U493 ( .A1(n681), .A2(n382), .ZN(n543) );
  NAND2_X1 U494 ( .A1(n531), .A2(n382), .ZN(n532) );
  NAND2_X1 U495 ( .A1(n594), .A2(n382), .ZN(n596) );
  NOR2_X1 U496 ( .A1(n569), .A2(n382), .ZN(n743) );
  AND2_X1 U497 ( .A1(n397), .A2(n347), .ZN(n652) );
  AND2_X1 U498 ( .A1(n641), .A2(G478), .ZN(n674) );
  NAND2_X1 U499 ( .A1(n454), .A2(G234), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n470), .A2(G221), .ZN(n439) );
  XNOR2_X2 U501 ( .A(n389), .B(n632), .ZN(n636) );
  NAND2_X1 U502 ( .A1(n635), .A2(KEYINPUT2), .ZN(n396) );
  INV_X1 U503 ( .A(KEYINPUT48), .ZN(n401) );
  INV_X1 U504 ( .A(KEYINPUT72), .ZN(n403) );
  NAND2_X1 U505 ( .A1(n404), .A2(n462), .ZN(n566) );
  XNOR2_X1 U506 ( .A(n406), .B(G119), .ZN(n415) );
  NAND2_X1 U507 ( .A1(n641), .A2(G210), .ZN(n667) );
  NAND2_X1 U508 ( .A1(n641), .A2(G472), .ZN(n658) );
  INV_X1 U509 ( .A(n519), .ZN(n571) );
  INV_X1 U510 ( .A(n745), .ZN(n407) );
  XNOR2_X1 U511 ( .A(n472), .B(n471), .ZN(n475) );
  INV_X1 U512 ( .A(n675), .ZN(n668) );
  NOR2_X1 U513 ( .A1(n454), .A2(G952), .ZN(n675) );
  XNOR2_X2 U514 ( .A(G128), .B(G143), .ZN(n501) );
  XNOR2_X1 U515 ( .A(KEYINPUT4), .B(G131), .ZN(n413) );
  NAND2_X1 U516 ( .A1(n483), .A2(G210), .ZN(n417) );
  XNOR2_X1 U517 ( .A(G137), .B(G101), .ZN(n416) );
  XNOR2_X1 U518 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U519 ( .A(KEYINPUT78), .B(KEYINPUT5), .ZN(n418) );
  XNOR2_X1 U520 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n495), .B(n420), .ZN(n421) );
  XNOR2_X1 U522 ( .A(n459), .B(n421), .ZN(n656) );
  XNOR2_X2 U523 ( .A(n422), .B(G472), .ZN(n563) );
  INV_X1 U524 ( .A(G902), .ZN(n488) );
  NAND2_X1 U525 ( .A1(n423), .A2(n488), .ZN(n508) );
  NAND2_X1 U526 ( .A1(n508), .A2(G214), .ZN(n424) );
  XNOR2_X1 U527 ( .A(n424), .B(KEYINPUT92), .ZN(n703) );
  XNOR2_X1 U528 ( .A(n425), .B(KEYINPUT30), .ZN(n431) );
  XNOR2_X1 U529 ( .A(KEYINPUT14), .B(n426), .ZN(n715) );
  NAND2_X1 U530 ( .A1(n488), .A2(G953), .ZN(n428) );
  AND2_X1 U531 ( .A1(n428), .A2(n427), .ZN(n429) );
  AND2_X1 U532 ( .A1(n715), .A2(n429), .ZN(n517) );
  NAND2_X1 U533 ( .A1(G953), .A2(G900), .ZN(n430) );
  AND2_X1 U534 ( .A1(n517), .A2(n430), .ZN(n526) );
  AND2_X1 U535 ( .A1(n431), .A2(n526), .ZN(n466) );
  XNOR2_X1 U536 ( .A(G110), .B(KEYINPUT24), .ZN(n434) );
  XNOR2_X1 U537 ( .A(n434), .B(n433), .ZN(n437) );
  XNOR2_X1 U538 ( .A(n435), .B(KEYINPUT75), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U540 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U541 ( .A(G146), .B(G125), .ZN(n503) );
  XNOR2_X1 U542 ( .A(n503), .B(KEYINPUT10), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G140), .B(G137), .ZN(n456) );
  XNOR2_X1 U544 ( .A(n485), .B(n456), .ZN(n584) );
  XNOR2_X1 U545 ( .A(n440), .B(n584), .ZN(n637) );
  NAND2_X1 U546 ( .A1(n633), .A2(G234), .ZN(n442) );
  XNOR2_X1 U547 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n442), .B(n441), .ZN(n447) );
  AND2_X1 U549 ( .A1(n447), .A2(G217), .ZN(n445) );
  XNOR2_X1 U550 ( .A(KEYINPUT80), .B(KEYINPUT95), .ZN(n443) );
  XNOR2_X1 U551 ( .A(n443), .B(KEYINPUT25), .ZN(n444) );
  XNOR2_X1 U552 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U553 ( .A1(n447), .A2(G221), .ZN(n449) );
  INV_X1 U554 ( .A(KEYINPUT21), .ZN(n448) );
  XNOR2_X1 U555 ( .A(n449), .B(n448), .ZN(n680) );
  INV_X1 U556 ( .A(n680), .ZN(n450) );
  XNOR2_X1 U557 ( .A(n451), .B(G110), .ZN(n453) );
  XNOR2_X1 U558 ( .A(G101), .B(KEYINPUT91), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n453), .B(n452), .ZN(n496) );
  NAND2_X1 U560 ( .A1(n454), .A2(G227), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U562 ( .A(n496), .B(n457), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n459), .B(n458), .ZN(n645) );
  XNOR2_X1 U564 ( .A(KEYINPUT73), .B(G469), .ZN(n460) );
  XNOR2_X2 U565 ( .A(n461), .B(n460), .ZN(n565) );
  INV_X1 U566 ( .A(n565), .ZN(n462) );
  NAND2_X1 U567 ( .A1(n546), .A2(n462), .ZN(n464) );
  INV_X1 U568 ( .A(KEYINPUT104), .ZN(n463) );
  XNOR2_X1 U569 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U570 ( .A1(n466), .A2(n465), .ZN(n467) );
  INV_X1 U571 ( .A(n557), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n470), .A2(G217), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n473), .B(G116), .ZN(n474) );
  XNOR2_X1 U574 ( .A(n475), .B(n474), .ZN(n672) );
  NAND2_X1 U575 ( .A1(n672), .A2(n488), .ZN(n476) );
  INV_X1 U576 ( .A(G478), .ZN(n671) );
  INV_X1 U577 ( .A(n554), .ZN(n492) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U579 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U580 ( .A(n482), .B(n481), .Z(n487) );
  AND2_X1 U581 ( .A1(n483), .A2(G214), .ZN(n484) );
  XNOR2_X1 U582 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U583 ( .A(n487), .B(n486), .ZN(n650) );
  NAND2_X1 U584 ( .A1(n650), .A2(n488), .ZN(n491) );
  XNOR2_X1 U585 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n489) );
  INV_X1 U586 ( .A(G475), .ZN(n649) );
  XNOR2_X1 U587 ( .A(n489), .B(n649), .ZN(n490) );
  XNOR2_X1 U588 ( .A(n491), .B(n490), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n492), .A2(n553), .ZN(n493) );
  XNOR2_X1 U590 ( .A(n493), .B(KEYINPUT101), .ZN(n605) );
  XNOR2_X1 U591 ( .A(n495), .B(n494), .ZN(n497) );
  XNOR2_X1 U592 ( .A(n497), .B(n496), .ZN(n751) );
  XNOR2_X1 U593 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n499) );
  NAND2_X1 U594 ( .A1(n454), .A2(G224), .ZN(n498) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U596 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U597 ( .A(KEYINPUT4), .B(KEYINPUT81), .ZN(n502) );
  XNOR2_X1 U598 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U599 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U600 ( .A(n751), .B(n506), .ZN(n664) );
  INV_X1 U601 ( .A(n664), .ZN(n507) );
  NAND2_X1 U602 ( .A1(n508), .A2(G210), .ZN(n510) );
  INV_X1 U603 ( .A(KEYINPUT83), .ZN(n509) );
  XNOR2_X1 U604 ( .A(n510), .B(n509), .ZN(n511) );
  BUF_X1 U605 ( .A(n515), .Z(n556) );
  INV_X1 U606 ( .A(n556), .ZN(n533) );
  NAND2_X1 U607 ( .A1(n605), .A2(n533), .ZN(n512) );
  NOR2_X1 U608 ( .A1(n513), .A2(n512), .ZN(n570) );
  XOR2_X1 U609 ( .A(G143), .B(n570), .Z(G45) );
  INV_X1 U610 ( .A(n703), .ZN(n514) );
  NAND2_X1 U611 ( .A1(G953), .A2(G898), .ZN(n516) );
  AND2_X1 U612 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n521), .B(n520), .ZN(n536) );
  NOR2_X1 U614 ( .A1(n691), .A2(n565), .ZN(n522) );
  NAND2_X1 U615 ( .A1(n522), .A2(n546), .ZN(n523) );
  OR2_X1 U616 ( .A1(n602), .A2(n523), .ZN(n727) );
  NOR2_X1 U617 ( .A1(n727), .A2(n551), .ZN(n524) );
  XOR2_X1 U618 ( .A(G104), .B(n524), .Z(G6) );
  XNOR2_X1 U619 ( .A(G140), .B(KEYINPUT112), .ZN(n535) );
  BUF_X1 U620 ( .A(n525), .Z(n597) );
  AND2_X1 U621 ( .A1(n680), .A2(n526), .ZN(n527) );
  XNOR2_X1 U622 ( .A(n563), .B(KEYINPUT6), .ZN(n608) );
  NAND2_X1 U623 ( .A1(n599), .A2(n738), .ZN(n528) );
  NAND2_X1 U624 ( .A1(n703), .A2(n568), .ZN(n529) );
  XNOR2_X1 U625 ( .A(n529), .B(KEYINPUT103), .ZN(n531) );
  XNOR2_X1 U626 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n530) );
  XOR2_X1 U627 ( .A(KEYINPUT43), .B(n532), .Z(n534) );
  NOR2_X1 U628 ( .A1(n534), .A2(n533), .ZN(n582) );
  XOR2_X1 U629 ( .A(n535), .B(n582), .Z(G42) );
  INV_X1 U630 ( .A(n536), .ZN(n538) );
  AND2_X1 U631 ( .A1(n554), .A2(n537), .ZN(n702) );
  XNOR2_X1 U632 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n540) );
  INV_X1 U633 ( .A(KEYINPUT65), .ZN(n539) );
  INV_X1 U634 ( .A(n610), .ZN(n594) );
  XNOR2_X1 U635 ( .A(n597), .B(KEYINPUT99), .ZN(n681) );
  NOR2_X1 U636 ( .A1(n543), .A2(n599), .ZN(n544) );
  NAND2_X1 U637 ( .A1(n594), .A2(n544), .ZN(n616) );
  XNOR2_X1 U638 ( .A(G101), .B(KEYINPUT110), .ZN(n545) );
  XNOR2_X1 U639 ( .A(n616), .B(n545), .ZN(G3) );
  INV_X1 U640 ( .A(n546), .ZN(n683) );
  XNOR2_X2 U641 ( .A(n547), .B(KEYINPUT77), .ZN(n690) );
  NAND2_X1 U642 ( .A1(n690), .A2(n691), .ZN(n548) );
  NOR2_X1 U643 ( .A1(n602), .A2(n548), .ZN(n550) );
  XNOR2_X1 U644 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n549) );
  XNOR2_X1 U645 ( .A(n550), .B(n549), .ZN(n614) );
  NOR2_X1 U646 ( .A1(n614), .A2(n551), .ZN(n552) );
  XOR2_X1 U647 ( .A(G113), .B(n552), .Z(G15) );
  OR2_X1 U648 ( .A1(n554), .A2(n553), .ZN(n732) );
  NOR2_X1 U649 ( .A1(n614), .A2(n732), .ZN(n555) );
  XOR2_X1 U650 ( .A(G116), .B(n555), .Z(G18) );
  XNOR2_X1 U651 ( .A(n556), .B(KEYINPUT38), .ZN(n704) );
  NAND2_X1 U652 ( .A1(n557), .A2(n704), .ZN(n559) );
  XNOR2_X1 U653 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n559), .B(n558), .ZN(n579) );
  NOR2_X2 U655 ( .A1(n579), .A2(n572), .ZN(n561) );
  XOR2_X1 U656 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n560) );
  XNOR2_X1 U657 ( .A(n561), .B(n560), .ZN(n662) );
  AND2_X1 U658 ( .A1(n704), .A2(n703), .ZN(n700) );
  NAND2_X1 U659 ( .A1(n700), .A2(n702), .ZN(n562) );
  INV_X1 U660 ( .A(n563), .ZN(n688) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT105), .ZN(n731) );
  NAND2_X1 U662 ( .A1(n719), .A2(n731), .ZN(n567) );
  XNOR2_X1 U663 ( .A(n567), .B(KEYINPUT42), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n743), .A2(n570), .ZN(n578) );
  NAND2_X1 U665 ( .A1(n572), .A2(n732), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n573), .B(KEYINPUT98), .ZN(n699) );
  NAND2_X1 U667 ( .A1(n699), .A2(KEYINPUT70), .ZN(n574) );
  NOR2_X1 U668 ( .A1(n571), .A2(n574), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n731), .A2(n575), .ZN(n576) );
  XOR2_X1 U670 ( .A(KEYINPUT47), .B(n576), .Z(n577) );
  OR2_X1 U671 ( .A1(n579), .A2(n732), .ZN(n581) );
  INV_X1 U672 ( .A(KEYINPUT108), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n581), .B(n580), .ZN(n758) );
  NOR2_X1 U674 ( .A1(n582), .A2(n758), .ZN(n583) );
  XNOR2_X1 U675 ( .A(n584), .B(KEYINPUT125), .ZN(n585) );
  XNOR2_X1 U676 ( .A(n586), .B(n585), .ZN(n588) );
  XNOR2_X1 U677 ( .A(n634), .B(n588), .ZN(n587) );
  NAND2_X1 U678 ( .A1(n587), .A2(n454), .ZN(n592) );
  XNOR2_X1 U679 ( .A(n588), .B(G227), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n589), .A2(G900), .ZN(n590) );
  NAND2_X1 U681 ( .A1(n590), .A2(G953), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n592), .A2(n591), .ZN(G72) );
  XNOR2_X1 U683 ( .A(n593), .B(G137), .ZN(G39) );
  INV_X1 U684 ( .A(n597), .ZN(n598) );
  XNOR2_X1 U685 ( .A(n622), .B(G110), .ZN(G12) );
  NAND2_X1 U686 ( .A1(n690), .A2(n599), .ZN(n601) );
  INV_X1 U687 ( .A(KEYINPUT33), .ZN(n600) );
  INV_X1 U688 ( .A(KEYINPUT34), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n604), .B(n603), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U691 ( .A(n607), .B(KEYINPUT35), .ZN(n670) );
  NAND2_X1 U692 ( .A1(n353), .A2(n608), .ZN(n609) );
  NOR2_X1 U693 ( .A1(n670), .A2(n613), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n614), .A2(n727), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n615), .A2(n699), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  INV_X1 U697 ( .A(n620), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n621), .A2(KEYINPUT44), .ZN(n624) );
  INV_X1 U699 ( .A(n622), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n670), .A2(KEYINPUT88), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n629) );
  INV_X1 U703 ( .A(KEYINPUT44), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n627), .A2(KEYINPUT88), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X1 U706 ( .A(KEYINPUT45), .ZN(n632) );
  INV_X1 U707 ( .A(n634), .ZN(n635) );
  BUF_X1 U708 ( .A(n636), .Z(n745) );
  NAND2_X1 U709 ( .A1(n641), .A2(G217), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT122), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n640), .A2(n675), .ZN(G66) );
  NAND2_X1 U713 ( .A1(n641), .A2(G469), .ZN(n647) );
  XOR2_X1 U714 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n643) );
  XNOR2_X1 U715 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n642) );
  XOR2_X1 U716 ( .A(n643), .B(n642), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n648), .A2(n675), .ZN(G54) );
  XOR2_X1 U720 ( .A(n650), .B(KEYINPUT59), .Z(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U722 ( .A1(n653), .A2(n675), .ZN(n655) );
  XNOR2_X1 U723 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G60) );
  XOR2_X1 U725 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n354), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n660) );
  XOR2_X1 U728 ( .A(G119), .B(KEYINPUT126), .Z(n661) );
  XNOR2_X1 U729 ( .A(n620), .B(n661), .ZN(G21) );
  XOR2_X1 U730 ( .A(G131), .B(KEYINPUT127), .Z(n663) );
  XNOR2_X1 U731 ( .A(n662), .B(n663), .ZN(G33) );
  BUF_X1 U732 ( .A(n664), .Z(n666) );
  XOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n665) );
  XNOR2_X1 U734 ( .A(n667), .B(n355), .ZN(n669) );
  XOR2_X1 U735 ( .A(G122), .B(n670), .Z(G24) );
  XOR2_X1 U736 ( .A(n672), .B(KEYINPUT121), .Z(n673) );
  XNOR2_X1 U737 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(G63) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n677) );
  NOR2_X1 U740 ( .A1(n410), .A2(n677), .ZN(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT84), .B(n678), .Z(n679) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U743 ( .A(n682), .B(KEYINPUT49), .ZN(n687) );
  XOR2_X1 U744 ( .A(KEYINPUT113), .B(KEYINPUT50), .Z(n684) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U746 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n694) );
  INV_X1 U748 ( .A(n690), .ZN(n692) );
  NAND2_X1 U749 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n695), .B(KEYINPUT114), .ZN(n696) );
  XOR2_X1 U752 ( .A(KEYINPUT51), .B(n696), .Z(n698) );
  INV_X1 U753 ( .A(n719), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n713) );
  NAND2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n701), .B(KEYINPUT117), .ZN(n710) );
  INV_X1 U757 ( .A(n702), .ZN(n707) );
  NOR2_X1 U758 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U759 ( .A(KEYINPUT115), .B(n705), .Z(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n708), .B(KEYINPUT116), .ZN(n709) );
  NOR2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n711), .A2(n718), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n714), .B(KEYINPUT52), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n715), .A2(G952), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n723) );
  NAND2_X1 U768 ( .A1(n381), .A2(n719), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n720), .B(KEYINPUT118), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n721), .A2(n454), .ZN(n722) );
  NOR2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U773 ( .A(KEYINPUT53), .B(n726), .Z(G75) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n729) );
  NOR2_X1 U775 ( .A1(n727), .A2(n732), .ZN(n728) );
  XOR2_X1 U776 ( .A(n729), .B(n728), .Z(n730) );
  XNOR2_X1 U777 ( .A(G107), .B(n730), .ZN(G9) );
  INV_X1 U778 ( .A(n731), .ZN(n741) );
  INV_X1 U779 ( .A(n571), .ZN(n739) );
  INV_X1 U780 ( .A(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n739), .A2(n733), .ZN(n734) );
  NOR2_X1 U782 ( .A1(n741), .A2(n734), .ZN(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT111), .B(KEYINPUT29), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n737) );
  XOR2_X1 U785 ( .A(G128), .B(n737), .Z(G30) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U787 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U788 ( .A(G146), .B(n742), .Z(G48) );
  XNOR2_X1 U789 ( .A(G125), .B(n743), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U791 ( .A1(n745), .A2(G953), .ZN(n750) );
  INV_X1 U792 ( .A(G898), .ZN(n748) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n746) );
  XOR2_X1 U794 ( .A(KEYINPUT61), .B(n746), .Z(n747) );
  NOR2_X1 U795 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U796 ( .A1(n750), .A2(n749), .ZN(n757) );
  BUF_X1 U797 ( .A(n751), .Z(n752) );
  XNOR2_X1 U798 ( .A(n752), .B(KEYINPUT123), .ZN(n754) );
  NOR2_X1 U799 ( .A1(n454), .A2(G898), .ZN(n753) );
  NOR2_X1 U800 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U801 ( .A(KEYINPUT124), .B(n755), .Z(n756) );
  XNOR2_X1 U802 ( .A(n757), .B(n756), .ZN(G69) );
  XOR2_X1 U803 ( .A(G134), .B(n758), .Z(G36) );
endmodule

