//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT2), .A2(G113), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G113), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT5), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n196), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G116), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT5), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n194), .A2(new_n199), .B1(new_n202), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n210), .A2(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n214), .B2(new_n217), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n206), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n196), .B2(new_n198), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n194), .ZN(new_n227));
  AND3_X1   g041(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(KEYINPUT2), .B2(G113), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT69), .B1(new_n203), .B2(new_n204), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n234), .A3(G101), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n221), .A2(new_n236), .A3(KEYINPUT82), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT82), .B1(new_n221), .B2(new_n236), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n224), .A2(new_n233), .A3(new_n235), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n194), .A2(new_n199), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n202), .A2(new_n205), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n214), .A2(new_n217), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT80), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n245), .B1(new_n246), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n221), .A2(new_n236), .A3(KEYINPUT82), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(new_n241), .A3(new_n243), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT84), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n259), .B(G146), .C1(new_n260), .C2(KEYINPUT1), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n266));
  OAI221_X1 g080(.A(new_n261), .B1(G128), .B2(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n263), .A2(new_n264), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n263), .A2(new_n264), .B1(KEYINPUT0), .B2(G128), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  OR2_X1    g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n268), .B1(new_n280), .B2(G125), .ZN(new_n281));
  INV_X1    g095(.A(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G224), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n281), .B(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n246), .A2(new_n253), .A3(new_n243), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n241), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n254), .A2(new_n243), .A3(new_n255), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n258), .B(new_n284), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n281), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n206), .A2(KEYINPUT85), .A3(new_n250), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n242), .B(KEYINPUT8), .ZN(new_n296));
  INV_X1    g110(.A(new_n250), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n249), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n206), .A2(KEYINPUT85), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n295), .B(new_n296), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n281), .A2(new_n293), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n294), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n285), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n294), .A2(KEYINPUT86), .A3(new_n301), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n291), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n291), .A2(new_n307), .A3(new_n309), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT87), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n291), .B2(new_n307), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n188), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT9), .B(G234), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G221), .B1(new_n319), .B2(G902), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT79), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G469), .ZN(new_n324));
  INV_X1    g138(.A(G902), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n297), .B(new_n267), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G131), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n332), .A3(new_n337), .A4(new_n333), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(KEYINPUT66), .A3(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT12), .B1(new_n327), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n267), .B(new_n250), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(new_n341), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n265), .A2(new_n277), .A3(new_n269), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT64), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(new_n274), .A3(new_n224), .A4(new_n235), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n297), .A2(new_n267), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT10), .B(new_n267), .C1(new_n219), .C2(new_n220), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .A4(new_n341), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n348), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G110), .B(G140), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n282), .A2(G227), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n363), .B(new_n364), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n358), .A2(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n358), .A2(new_n359), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n342), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n362), .A2(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n326), .B1(new_n372), .B2(G469), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n348), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n371), .B1(new_n360), .B2(new_n361), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n366), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n324), .A3(new_n325), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n323), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G478), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(KEYINPUT15), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n319), .A2(new_n382), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n260), .B2(G143), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT90), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n259), .A2(G128), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n389), .B(new_n384), .C1(new_n260), .C2(G143), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n260), .A2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n386), .A2(KEYINPUT91), .A3(new_n388), .A4(new_n390), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G134), .ZN(new_n398));
  INV_X1    g212(.A(G122), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT89), .B1(new_n399), .B2(G116), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n195), .A3(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n195), .B2(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G107), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n403), .B(new_n210), .C1(new_n195), .C2(G122), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n394), .A2(new_n387), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n405), .A2(new_n406), .B1(new_n329), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT92), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n407), .B(new_n329), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n415), .A2(KEYINPUT93), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(KEYINPUT93), .ZN(new_n417));
  OAI22_X1  g231(.A1(new_n403), .A2(KEYINPUT14), .B1(new_n195), .B2(G122), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n406), .B(new_n414), .C1(new_n419), .C2(new_n210), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n383), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n398), .A2(new_n411), .A3(new_n408), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n411), .B1(new_n398), .B2(new_n408), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n420), .B(new_n383), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n325), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n381), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  INV_X1    g244(.A(new_n383), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(G902), .B1(new_n432), .B2(new_n424), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT94), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n428), .B1(new_n435), .B2(new_n381), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n282), .A3(G214), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n259), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G131), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(G143), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n337), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT17), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(G125), .ZN(new_n449));
  INV_X1    g263(.A(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G140), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n448), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(G146), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n445), .B(new_n454), .C1(new_n444), .C2(new_n441), .ZN(new_n455));
  XNOR2_X1  g269(.A(G113), .B(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(new_n207), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT18), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n442), .B1(new_n458), .B2(new_n337), .ZN(new_n459));
  XNOR2_X1  g273(.A(G125), .B(G140), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(new_n262), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n459), .B(new_n461), .C1(new_n458), .C2(new_n441), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n460), .B(KEYINPUT19), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n262), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n453), .A2(new_n262), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n442), .A2(new_n337), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n440), .A2(G131), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n462), .ZN(new_n470));
  INV_X1    g284(.A(new_n457), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n463), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n463), .B2(new_n472), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT20), .B(new_n437), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n472), .ZN(new_n477));
  INV_X1    g291(.A(new_n463), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n437), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n457), .B1(new_n455), .B2(new_n462), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n325), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G475), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n282), .A2(G952), .ZN(new_n486));
  NAND2_X1  g300(.A1(G234), .A2(G237), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(G902), .A3(G953), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n379), .A2(new_n436), .A3(new_n485), .A4(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n187), .B1(new_n317), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n188), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n291), .A2(new_n307), .A3(new_n309), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n315), .B1(new_n495), .B2(new_n314), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n311), .A2(KEYINPUT87), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n432), .A2(new_n424), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT94), .B1(new_n499), .B2(new_n325), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n427), .B(G902), .C1(new_n432), .C2(new_n424), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n381), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n433), .A2(KEYINPUT94), .B1(KEYINPUT15), .B2(new_n380), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(new_n505));
  INV_X1    g319(.A(new_n491), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n498), .A2(KEYINPUT95), .A3(new_n379), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n280), .B2(new_n341), .ZN(new_n511));
  INV_X1    g325(.A(new_n333), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n329), .A2(G137), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n267), .A2(new_n338), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n350), .A2(new_n351), .B1(new_n270), .B2(new_n273), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(KEYINPUT67), .A3(new_n340), .A4(new_n339), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n352), .A2(new_n340), .A3(new_n339), .A4(new_n274), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n521), .A2(KEYINPUT30), .A3(new_n515), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n233), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n515), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n233), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n438), .A2(new_n282), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n212), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n524), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n522), .B1(new_n518), .B2(new_n519), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n526), .B1(new_n536), .B2(new_n233), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n532), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n227), .B(new_n232), .C1(new_n525), .C2(KEYINPUT71), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n521), .B2(new_n515), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n526), .B1(new_n233), .B2(new_n518), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(new_n539), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n535), .A2(new_n538), .B1(new_n545), .B2(new_n531), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n509), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n531), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n533), .A2(new_n534), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT31), .B1(new_n537), .B2(new_n532), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n547), .ZN(new_n554));
  INV_X1    g368(.A(new_n531), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n531), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT29), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n525), .B(new_n233), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n543), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n325), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G472), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n549), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n382), .B1(G234), .B2(new_n325), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n568));
  XNOR2_X1  g382(.A(G119), .B(G128), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT72), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT24), .B(G110), .Z(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT73), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT74), .B1(new_n197), .B2(G128), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n575), .A2(KEYINPUT23), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n197), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(KEYINPUT23), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n454), .B1(G110), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT72), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n569), .B(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n584), .B2(new_n571), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT75), .B(G110), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n570), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  MUX2_X1   g404(.A(new_n452), .B(new_n453), .S(G146), .Z(new_n591));
  AND3_X1   g405(.A1(new_n590), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT77), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n581), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n282), .A2(G221), .A3(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n581), .B(new_n597), .C1(new_n592), .C2(new_n593), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n568), .B1(new_n601), .B2(G902), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n599), .A2(KEYINPUT25), .A3(new_n325), .A4(new_n600), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n567), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n601), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n566), .A2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n565), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n493), .A2(new_n508), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  NAND2_X1  g426(.A1(new_n553), .A2(new_n325), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n613), .A2(G472), .B1(new_n553), .B2(new_n547), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n614), .A2(new_n609), .A3(new_n379), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n494), .B1(new_n311), .B2(new_n312), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n491), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n432), .A2(KEYINPUT33), .A3(new_n424), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT33), .B1(new_n432), .B2(new_n424), .ZN(new_n622));
  OAI21_X1  g436(.A(G478), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n433), .A2(new_n380), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n380), .A2(new_n325), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n623), .A2(new_n505), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  NAND2_X1  g445(.A1(new_n476), .A2(new_n484), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n474), .A2(new_n475), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT20), .B1(new_n633), .B2(new_n437), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n436), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT96), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(new_n604), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n594), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n606), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n493), .A2(new_n508), .A3(new_n614), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n488), .B(KEYINPUT97), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  INV_X1    g464(.A(new_n490), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n634), .A2(new_n632), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n648), .B1(new_n504), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n504), .A2(new_n648), .A3(new_n653), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n565), .A2(new_n379), .A3(new_n616), .A4(new_n644), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n260), .ZN(G30));
  NOR2_X1   g474(.A1(new_n313), .A2(new_n316), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT38), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n652), .B(KEYINPUT39), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n379), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n604), .B1(new_n642), .B2(new_n606), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n665), .B2(KEYINPUT40), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n537), .A2(new_n531), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n325), .B1(new_n559), .B2(new_n555), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n549), .A2(new_n554), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(new_n188), .A3(new_n504), .A4(new_n505), .ZN(new_n673));
  OR4_X1    g487(.A1(new_n662), .A2(new_n666), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  NOR2_X1   g489(.A1(new_n627), .A2(new_n652), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n658), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n262), .ZN(G48));
  AOI22_X1  g493(.A1(new_n348), .A2(new_n369), .B1(new_n375), .B2(new_n366), .ZN(new_n680));
  OAI21_X1  g494(.A(G469), .B1(new_n680), .B2(G902), .ZN(new_n681));
  INV_X1    g495(.A(new_n321), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n378), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT99), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n378), .A3(new_n685), .A4(new_n682), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n610), .A2(new_n628), .A3(new_n618), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  AND3_X1   g504(.A1(new_n684), .A2(new_n616), .A3(new_n686), .ZN(new_n691));
  INV_X1    g505(.A(new_n609), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n506), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n693), .A3(new_n565), .A4(new_n635), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT100), .B(G116), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G18));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n565), .A3(new_n507), .A4(new_n644), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  AND4_X1   g512(.A1(new_n491), .A2(new_n684), .A3(new_n616), .A4(new_n686), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n604), .A2(new_n608), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n535), .A2(new_n538), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n550), .ZN(new_n706));
  INV_X1    g520(.A(G472), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(KEYINPUT102), .B(G472), .C1(new_n546), .C2(G902), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n561), .A2(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n561), .A2(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n531), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n708), .A2(new_n709), .B1(new_n547), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n436), .B2(new_n485), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n504), .A2(KEYINPUT104), .A3(new_n505), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n699), .A2(new_n703), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n547), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT102), .B1(new_n613), .B2(G472), .ZN(new_n722));
  INV_X1    g536(.A(new_n709), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n644), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n676), .A2(new_n684), .A3(new_n616), .A4(new_n686), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n450), .ZN(G27));
  AOI21_X1  g541(.A(new_n321), .B1(new_n373), .B2(new_n378), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n676), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n496), .A2(new_n188), .A3(new_n497), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n610), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n731), .A2(new_n735), .A3(new_n610), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n549), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT106), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n553), .A2(new_n547), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT106), .A3(new_n509), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n554), .A3(new_n564), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n703), .A4(new_n731), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  INV_X1    g559(.A(new_n565), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n730), .A3(new_n692), .ZN(new_n747));
  INV_X1    g561(.A(new_n656), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT107), .B1(new_n748), .B2(new_n654), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n655), .A2(new_n750), .A3(new_n656), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n747), .A2(new_n749), .A3(new_n728), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  INV_X1    g567(.A(new_n622), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n620), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n625), .B1(new_n755), .B2(G478), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n624), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n757), .B2(new_n505), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n759), .A3(new_n485), .A4(new_n624), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n614), .A2(new_n667), .A3(KEYINPUT109), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT109), .B1(new_n614), .B2(new_n667), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n730), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT108), .Z(new_n773));
  INV_X1    g587(.A(new_n326), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n378), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n682), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n769), .A2(new_n663), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n331), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n682), .C1(new_n776), .C2(new_n777), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n677), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n730), .A2(new_n565), .A3(new_n609), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n719), .A2(new_n688), .A3(new_n694), .A4(new_n697), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n744), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n789), .B1(new_n792), .B2(KEYINPUT115), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n188), .B(new_n491), .C1(new_n313), .C2(new_n316), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT110), .B1(new_n794), .B2(new_n627), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n498), .A2(new_n628), .A3(new_n796), .A4(new_n491), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n615), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n504), .A2(new_n485), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT111), .ZN(new_n800));
  INV_X1    g614(.A(new_n794), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n615), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n645), .A3(new_n611), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n708), .A2(new_n709), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n680), .A2(G469), .A3(G902), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n371), .B(new_n365), .C1(new_n360), .C2(new_n361), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n347), .B1(new_n367), .B2(new_n368), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n365), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n324), .B1(new_n808), .B2(new_n325), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n682), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n627), .A3(new_n652), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n811), .A3(new_n721), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n565), .A2(new_n379), .A3(new_n436), .A4(new_n653), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n644), .A3(new_n767), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n752), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n803), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n658), .B1(new_n657), .B2(new_n677), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n726), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT104), .B1(new_n504), .B2(new_n505), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n715), .B(new_n485), .C1(new_n502), .C2(new_n503), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n616), .B(new_n672), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n652), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n667), .A2(new_n823), .A3(new_n728), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT112), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n188), .B1(new_n495), .B2(new_n314), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n716), .B2(new_n717), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n644), .A2(new_n652), .A3(new_n810), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n672), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n819), .A2(new_n831), .A3(KEYINPUT52), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n819), .B2(new_n831), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n790), .B1(new_n737), .B2(new_n743), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n793), .A2(new_n817), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n817), .B(new_n835), .C1(new_n833), .C2(new_n832), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n839), .B2(new_n842), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n788), .B(new_n838), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n839), .B2(new_n841), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n788), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n703), .A2(new_n714), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n649), .A3(new_n761), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n691), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n681), .A2(new_n378), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n782), .B(new_n783), .C1(new_n322), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n767), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n767), .A2(new_n687), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n860), .A2(new_n692), .A3(new_n488), .A4(new_n672), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n485), .A3(new_n757), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n761), .A2(new_n649), .A3(new_n687), .A4(new_n767), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n724), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n662), .A2(new_n494), .A3(new_n687), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(KEYINPUT50), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n859), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n742), .A2(new_n703), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n872), .A2(new_n863), .A3(KEYINPUT117), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT117), .B1(new_n872), .B2(new_n863), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT48), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n486), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n861), .A2(new_n628), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n870), .A3(KEYINPUT51), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n856), .A2(new_n881), .B1(G952), .B2(G953), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n188), .A3(new_n322), .A4(new_n884), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n885), .A2(new_n672), .A3(new_n700), .A4(new_n702), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n757), .A2(new_n505), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n662), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n882), .A2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n282), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(G210), .A3(G902), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n258), .B1(new_n289), .B2(new_n290), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n284), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n893), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n894), .B1(new_n893), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n892), .A2(KEYINPUT118), .A3(G210), .A4(G902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n898), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n897), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n902), .A2(new_n907), .ZN(G51));
  NAND2_X1  g722(.A1(new_n774), .A2(KEYINPUT57), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n774), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n839), .A2(new_n842), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT114), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n788), .B1(new_n914), .B2(new_n838), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n909), .B(new_n910), .C1(new_n915), .C2(new_n846), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n377), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n325), .B1(new_n914), .B2(new_n838), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n773), .B(KEYINPUT120), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n890), .B1(new_n917), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n633), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n890), .ZN(G60));
  XNOR2_X1  g740(.A(new_n625), .B(KEYINPUT59), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n755), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n915), .B2(new_n846), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n891), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n845), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n934), .B2(new_n890), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n755), .B1(new_n850), .B2(new_n927), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n930), .A2(new_n935), .A3(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n892), .A2(new_n642), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n891), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n605), .B1(new_n892), .B2(new_n939), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n943), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n940), .A2(new_n891), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n944), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n946), .A2(new_n950), .ZN(G66));
  NOR2_X1   g765(.A1(new_n803), .A2(new_n790), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(G953), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n489), .A2(G224), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n282), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n895), .B1(G898), .B2(new_n282), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  XNOR2_X1  g772(.A(new_n536), .B(KEYINPUT124), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n464), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n819), .A2(new_n752), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n784), .B2(new_n785), .ZN(new_n962));
  INV_X1    g776(.A(new_n827), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n769), .B1(new_n872), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n778), .A2(new_n663), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n964), .A2(new_n965), .B1(new_n737), .B2(new_n743), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n282), .A2(G900), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT125), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n968), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n960), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G227), .A2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(G953), .ZN(new_n974));
  INV_X1    g788(.A(new_n960), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n800), .A2(new_n628), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n665), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n779), .B1(new_n747), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n674), .A2(new_n819), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT62), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n980), .A3(new_n786), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n975), .B1(new_n982), .B2(G953), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n972), .A2(new_n974), .A3(new_n983), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n968), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n969), .ZN(new_n986));
  OAI211_X1 g800(.A(G953), .B(new_n973), .C1(new_n986), .C2(new_n975), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G72));
  NAND3_X1  g802(.A1(new_n962), .A2(new_n952), .A3(new_n966), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n557), .B1(new_n992), .B2(KEYINPUT127), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n890), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n848), .ZN(new_n996));
  INV_X1    g810(.A(new_n669), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n557), .A3(new_n997), .A4(new_n991), .ZN(new_n998));
  INV_X1    g812(.A(new_n952), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n991), .B1(new_n981), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1002), .B(new_n991), .C1(new_n981), .C2(new_n999), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1001), .A2(new_n669), .A3(new_n1003), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n995), .A2(new_n998), .A3(new_n1004), .ZN(G57));
endmodule


