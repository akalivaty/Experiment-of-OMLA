

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729;

  NOR2_X1 U377 ( .A1(n522), .A2(n533), .ZN(n661) );
  INV_X1 U378 ( .A(G953), .ZN(n448) );
  NOR2_X1 U379 ( .A1(n644), .A2(n511), .ZN(n615) );
  AND2_X4 U380 ( .A1(n423), .A2(n637), .ZN(n697) );
  NOR2_X2 U381 ( .A1(n531), .A2(n409), .ZN(n408) );
  XNOR2_X2 U382 ( .A(n442), .B(n441), .ZN(n644) );
  XNOR2_X1 U383 ( .A(n519), .B(KEYINPUT66), .ZN(n641) );
  INV_X1 U384 ( .A(G113), .ZN(n406) );
  INV_X4 U385 ( .A(G131), .ZN(n443) );
  XNOR2_X1 U386 ( .A(n408), .B(n359), .ZN(n513) );
  AND2_X1 U387 ( .A1(n529), .A2(n578), .ZN(n520) );
  XNOR2_X1 U388 ( .A(n556), .B(n425), .ZN(n595) );
  INV_X1 U389 ( .A(n641), .ZN(n355) );
  XNOR2_X1 U390 ( .A(n707), .B(KEYINPUT74), .ZN(n482) );
  XNOR2_X1 U391 ( .A(n405), .B(n480), .ZN(n510) );
  XNOR2_X1 U392 ( .A(n454), .B(n453), .ZN(n707) );
  XNOR2_X1 U393 ( .A(n445), .B(G134), .ZN(n463) );
  XNOR2_X1 U394 ( .A(n483), .B(n391), .ZN(n714) );
  XNOR2_X1 U395 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U396 ( .A(n444), .B(KEYINPUT70), .ZN(n383) );
  INV_X1 U397 ( .A(G137), .ZN(n444) );
  XNOR2_X1 U398 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n432) );
  XOR2_X1 U399 ( .A(G107), .B(G104), .Z(n453) );
  XNOR2_X1 U400 ( .A(KEYINPUT92), .B(G101), .ZN(n452) );
  XNOR2_X1 U401 ( .A(G119), .B(G116), .ZN(n407) );
  XNOR2_X2 U402 ( .A(n403), .B(n357), .ZN(n596) );
  XNOR2_X1 U403 ( .A(n463), .B(n381), .ZN(n509) );
  XNOR2_X1 U404 ( .A(n446), .B(n382), .ZN(n381) );
  XNOR2_X1 U405 ( .A(n473), .B(n383), .ZN(n382) );
  INV_X1 U406 ( .A(KEYINPUT81), .ZN(n419) );
  XNOR2_X1 U407 ( .A(n398), .B(n396), .ZN(n458) );
  XNOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n398) );
  NOR2_X1 U409 ( .A1(n397), .A2(G953), .ZN(n396) );
  INV_X1 U410 ( .A(G234), .ZN(n397) );
  XOR2_X1 U411 ( .A(G125), .B(G146), .Z(n483) );
  AND2_X1 U412 ( .A1(n595), .A2(n355), .ZN(n529) );
  INV_X1 U413 ( .A(n595), .ZN(n640) );
  INV_X1 U414 ( .A(KEYINPUT88), .ZN(n599) );
  OR2_X2 U415 ( .A1(n605), .A2(G902), .ZN(n415) );
  XNOR2_X1 U416 ( .A(n465), .B(n464), .ZN(n692) );
  XNOR2_X1 U417 ( .A(G107), .B(G122), .ZN(n462) );
  XNOR2_X1 U418 ( .A(n713), .B(n372), .ZN(n680) );
  XNOR2_X1 U419 ( .A(n482), .B(n373), .ZN(n372) );
  XNOR2_X1 U420 ( .A(n451), .B(n455), .ZN(n373) );
  XNOR2_X1 U421 ( .A(n400), .B(KEYINPUT41), .ZN(n655) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n425) );
  XNOR2_X1 U423 ( .A(n585), .B(n492), .ZN(n558) );
  XNOR2_X1 U424 ( .A(n509), .B(n416), .ZN(n605) );
  XNOR2_X1 U425 ( .A(n436), .B(n390), .ZN(n698) );
  XNOR2_X1 U426 ( .A(n356), .B(n714), .ZN(n390) );
  NAND2_X1 U427 ( .A1(n421), .A2(n420), .ZN(n423) );
  NAND2_X1 U428 ( .A1(n424), .A2(KEYINPUT2), .ZN(n420) );
  NAND2_X1 U429 ( .A1(n697), .A2(G210), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n379), .B(n404), .ZN(n378) );
  INV_X1 U431 ( .A(KEYINPUT87), .ZN(n404) );
  AND2_X1 U432 ( .A1(n634), .A2(n597), .ZN(n601) );
  XOR2_X1 U433 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n460) );
  XNOR2_X1 U434 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  XNOR2_X1 U435 ( .A(n589), .B(KEYINPUT89), .ZN(n590) );
  AND2_X1 U436 ( .A1(n601), .A2(KEYINPUT2), .ZN(n598) );
  XNOR2_X1 U437 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U438 ( .A(n484), .B(n427), .ZN(n485) );
  XNOR2_X1 U439 ( .A(n445), .B(n483), .ZN(n486) );
  AND2_X1 U440 ( .A1(G224), .A2(n448), .ZN(n427) );
  NAND2_X1 U441 ( .A1(G237), .A2(G234), .ZN(n493) );
  NOR2_X1 U442 ( .A1(n571), .A2(n658), .ZN(n664) );
  NAND2_X1 U443 ( .A1(n661), .A2(n643), .ZN(n409) );
  INV_X1 U444 ( .A(n552), .ZN(n374) );
  XNOR2_X1 U445 ( .A(G146), .B(G101), .ZN(n504) );
  XOR2_X1 U446 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n505) );
  AND2_X1 U447 ( .A1(n602), .A2(n601), .ZN(n719) );
  XNOR2_X1 U448 ( .A(G122), .B(KEYINPUT16), .ZN(n481) );
  XNOR2_X1 U449 ( .A(G128), .B(G110), .ZN(n430) );
  XNOR2_X1 U450 ( .A(G122), .B(G113), .ZN(n467) );
  XNOR2_X1 U451 ( .A(KEYINPUT10), .B(G140), .ZN(n391) );
  AND2_X1 U452 ( .A1(n719), .A2(n424), .ZN(n365) );
  INV_X1 U453 ( .A(n603), .ZN(n424) );
  AND2_X1 U454 ( .A1(n638), .A2(n637), .ZN(n380) );
  NOR2_X1 U455 ( .A1(n701), .A2(KEYINPUT2), .ZN(n636) );
  NOR2_X1 U456 ( .A1(n580), .A2(n579), .ZN(n581) );
  AND2_X1 U457 ( .A1(n595), .A2(n370), .ZN(n512) );
  INV_X1 U458 ( .A(n644), .ZN(n370) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n534) );
  XNOR2_X1 U460 ( .A(n466), .B(G478), .ZN(n401) );
  OR2_X1 U461 ( .A1(n692), .A2(G902), .ZN(n402) );
  NOR2_X1 U462 ( .A1(G902), .A2(n680), .ZN(n457) );
  INV_X1 U463 ( .A(KEYINPUT0), .ZN(n410) );
  XOR2_X1 U464 ( .A(n546), .B(KEYINPUT6), .Z(n578) );
  AND2_X1 U465 ( .A1(n412), .A2(n548), .ZN(n635) );
  XNOR2_X1 U466 ( .A(n413), .B(KEYINPUT43), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n584), .A2(n414), .ZN(n413) );
  NOR2_X1 U468 ( .A1(n595), .A2(n663), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n573), .B(KEYINPUT42), .ZN(n727) );
  NAND2_X1 U470 ( .A1(n388), .A2(n392), .ZN(n387) );
  XNOR2_X1 U471 ( .A(n389), .B(n361), .ZN(n388) );
  AND2_X1 U472 ( .A1(n393), .A2(n392), .ZN(n700) );
  XNOR2_X1 U473 ( .A(n395), .B(n394), .ZN(n393) );
  INV_X1 U474 ( .A(n698), .ZN(n394) );
  INV_X1 U475 ( .A(KEYINPUT123), .ZN(n411) );
  INV_X1 U476 ( .A(KEYINPUT56), .ZN(n366) );
  NAND2_X1 U477 ( .A1(n368), .A2(n392), .ZN(n367) );
  XNOR2_X1 U478 ( .A(n369), .B(n360), .ZN(n368) );
  NAND2_X1 U479 ( .A1(n378), .A2(n429), .ZN(n363) );
  XOR2_X1 U480 ( .A(n431), .B(n430), .Z(n356) );
  AND2_X1 U481 ( .A1(G210), .A2(n491), .ZN(n357) );
  XNOR2_X1 U482 ( .A(n457), .B(n456), .ZN(n556) );
  XOR2_X1 U483 ( .A(n639), .B(KEYINPUT86), .Z(n358) );
  XNOR2_X1 U484 ( .A(n509), .B(n447), .ZN(n713) );
  XOR2_X1 U485 ( .A(n503), .B(KEYINPUT64), .Z(n359) );
  XOR2_X1 U486 ( .A(n679), .B(n426), .Z(n360) );
  XOR2_X1 U487 ( .A(n605), .B(n604), .Z(n361) );
  NOR2_X1 U488 ( .A1(G952), .A2(n448), .ZN(n699) );
  INV_X1 U489 ( .A(n699), .ZN(n392) );
  NAND2_X1 U490 ( .A1(n362), .A2(n554), .ZN(n511) );
  INV_X1 U491 ( .A(n537), .ZN(n362) );
  XNOR2_X1 U492 ( .A(n363), .B(n678), .ZN(G75) );
  NAND2_X1 U493 ( .A1(n364), .A2(n724), .ZN(n418) );
  XNOR2_X1 U494 ( .A(n518), .B(n517), .ZN(n364) );
  NAND2_X1 U495 ( .A1(n513), .A2(n514), .ZN(n515) );
  NAND2_X1 U496 ( .A1(n417), .A2(n541), .ZN(n542) );
  NOR2_X2 U497 ( .A1(n695), .A2(n699), .ZN(n696) );
  NAND2_X1 U498 ( .A1(n701), .A2(n365), .ZN(n421) );
  XNOR2_X2 U499 ( .A(n542), .B(KEYINPUT45), .ZN(n701) );
  XNOR2_X1 U500 ( .A(n367), .B(n366), .ZN(G51) );
  XNOR2_X2 U501 ( .A(n371), .B(n419), .ZN(n445) );
  XNOR2_X2 U502 ( .A(G128), .B(G143), .ZN(n371) );
  AND2_X1 U503 ( .A1(n375), .A2(n374), .ZN(n547) );
  XNOR2_X1 U504 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U505 ( .A(KEYINPUT30), .ZN(n376) );
  NAND2_X1 U506 ( .A1(n546), .A2(n593), .ZN(n377) );
  XNOR2_X2 U507 ( .A(n415), .B(G472), .ZN(n546) );
  NAND2_X1 U508 ( .A1(n380), .A2(n358), .ZN(n379) );
  NOR2_X1 U509 ( .A1(n641), .A2(n556), .ZN(n386) );
  NAND2_X1 U510 ( .A1(n384), .A2(n355), .ZN(n566) );
  AND2_X1 U511 ( .A1(n547), .A2(n385), .ZN(n384) );
  INV_X1 U512 ( .A(n556), .ZN(n385) );
  NAND2_X1 U513 ( .A1(n532), .A2(n386), .ZN(n609) );
  XNOR2_X1 U514 ( .A(n387), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U515 ( .A1(n697), .A2(G472), .ZN(n389) );
  NAND2_X1 U516 ( .A1(n697), .A2(G217), .ZN(n395) );
  INV_X1 U517 ( .A(n655), .ZN(n673) );
  NAND2_X1 U518 ( .A1(n655), .A2(n399), .ZN(n573) );
  INV_X1 U519 ( .A(n572), .ZN(n399) );
  NAND2_X1 U520 ( .A1(n664), .A2(n593), .ZN(n400) );
  NOR2_X2 U521 ( .A1(n551), .A2(n550), .ZN(n622) );
  NAND2_X1 U522 ( .A1(n596), .A2(n593), .ZN(n585) );
  NAND2_X1 U523 ( .A1(n679), .A2(n603), .ZN(n403) );
  XNOR2_X2 U524 ( .A(n500), .B(n410), .ZN(n531) );
  XNOR2_X1 U525 ( .A(n696), .B(n411), .ZN(G63) );
  XNOR2_X1 U526 ( .A(n510), .B(n508), .ZN(n416) );
  NAND2_X1 U527 ( .A1(n418), .A2(n528), .ZN(n417) );
  INV_X1 U528 ( .A(n526), .ZN(n724) );
  XNOR2_X1 U529 ( .A(n600), .B(n599), .ZN(n422) );
  NAND2_X1 U530 ( .A1(n422), .A2(n701), .ZN(n637) );
  NOR2_X2 U531 ( .A1(n690), .A2(n699), .ZN(n691) );
  XNOR2_X1 U532 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U533 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n426) );
  AND2_X1 U534 ( .A1(n506), .A2(G210), .ZN(n428) );
  NOR2_X1 U535 ( .A1(n677), .A2(G953), .ZN(n429) );
  INV_X1 U536 ( .A(KEYINPUT79), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n507), .B(n428), .ZN(n508) );
  XNOR2_X1 U538 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U539 ( .A(n452), .B(G110), .ZN(n454) );
  XNOR2_X1 U540 ( .A(n591), .B(n590), .ZN(n602) );
  XNOR2_X1 U541 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U542 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U543 ( .A(n689), .B(n688), .ZN(n690) );
  INV_X1 U544 ( .A(n727), .ZN(n728) );
  XOR2_X1 U545 ( .A(G137), .B(G119), .Z(n431) );
  XNOR2_X1 U546 ( .A(n432), .B(KEYINPUT23), .ZN(n433) );
  XOR2_X1 U547 ( .A(KEYINPUT96), .B(n433), .Z(n435) );
  NAND2_X1 U548 ( .A1(G221), .A2(n458), .ZN(n434) );
  XNOR2_X1 U549 ( .A(n435), .B(n434), .ZN(n436) );
  NOR2_X1 U550 ( .A1(G902), .A2(n698), .ZN(n442) );
  XOR2_X1 U551 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n439) );
  NAND2_X1 U552 ( .A1(G234), .A2(n603), .ZN(n437) );
  XNOR2_X1 U553 ( .A(KEYINPUT20), .B(n437), .ZN(n501) );
  NAND2_X1 U554 ( .A1(n501), .A2(G217), .ZN(n438) );
  XNOR2_X1 U555 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U556 ( .A(KEYINPUT97), .B(n440), .ZN(n441) );
  INV_X1 U557 ( .A(KEYINPUT95), .ZN(n447) );
  XNOR2_X2 U558 ( .A(n443), .B(KEYINPUT69), .ZN(n473) );
  XOR2_X1 U559 ( .A(KEYINPUT4), .B(KEYINPUT67), .Z(n484) );
  INV_X1 U560 ( .A(n484), .ZN(n446) );
  NAND2_X1 U561 ( .A1(G227), .A2(n448), .ZN(n450) );
  XNOR2_X1 U562 ( .A(G146), .B(G140), .ZN(n455) );
  XNOR2_X1 U563 ( .A(KEYINPUT72), .B(G469), .ZN(n456) );
  NAND2_X1 U564 ( .A1(G217), .A2(n458), .ZN(n459) );
  XNOR2_X1 U565 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U566 ( .A(n461), .B(G116), .Z(n465) );
  XNOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n466) );
  INV_X1 U568 ( .A(n534), .ZN(n522) );
  XOR2_X1 U569 ( .A(KEYINPUT99), .B(G143), .Z(n468) );
  XNOR2_X1 U570 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U571 ( .A(n714), .B(n469), .ZN(n477) );
  XOR2_X1 U572 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n471) );
  NOR2_X1 U573 ( .A1(G953), .A2(G237), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n506), .A2(G214), .ZN(n470) );
  XNOR2_X1 U575 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U576 ( .A(G104), .B(n472), .ZN(n475) );
  INV_X1 U577 ( .A(n473), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n687) );
  NOR2_X1 U580 ( .A1(G902), .A2(n687), .ZN(n479) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(G475), .ZN(n478) );
  XNOR2_X1 U582 ( .A(n479), .B(n478), .ZN(n533) );
  XNOR2_X1 U583 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n492) );
  XNOR2_X1 U584 ( .A(KEYINPUT3), .B(KEYINPUT73), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n481), .B(n510), .ZN(n706) );
  XNOR2_X1 U586 ( .A(n482), .B(n706), .ZN(n490) );
  XNOR2_X1 U587 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n487) );
  XNOR2_X1 U588 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n490), .B(n489), .ZN(n679) );
  OR2_X1 U590 ( .A1(G902), .A2(G237), .ZN(n491) );
  NAND2_X1 U591 ( .A1(G214), .A2(n491), .ZN(n593) );
  XOR2_X1 U592 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n494) );
  XNOR2_X1 U593 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U594 ( .A1(G952), .A2(n495), .ZN(n671) );
  NOR2_X1 U595 ( .A1(G953), .A2(n671), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G902), .A2(n495), .ZN(n496) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(n496), .Z(n497) );
  NAND2_X1 U598 ( .A1(G953), .A2(n497), .ZN(n543) );
  NOR2_X1 U599 ( .A1(G898), .A2(n543), .ZN(n498) );
  NOR2_X1 U600 ( .A1(n545), .A2(n498), .ZN(n499) );
  NOR2_X2 U601 ( .A1(n558), .A2(n499), .ZN(n500) );
  NAND2_X1 U602 ( .A1(n501), .A2(G221), .ZN(n502) );
  XOR2_X1 U603 ( .A(KEYINPUT21), .B(n502), .Z(n643) );
  XOR2_X1 U604 ( .A(KEYINPUT22), .B(KEYINPUT76), .Z(n503) );
  NAND2_X1 U605 ( .A1(n640), .A2(n513), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n505), .B(n504), .ZN(n507) );
  INV_X1 U607 ( .A(n546), .ZN(n554) );
  XNOR2_X1 U608 ( .A(n512), .B(KEYINPUT104), .ZN(n514) );
  NOR2_X1 U609 ( .A1(n515), .A2(n578), .ZN(n516) );
  XNOR2_X1 U610 ( .A(n516), .B(KEYINPUT32), .ZN(n726) );
  NOR2_X1 U611 ( .A1(n615), .A2(n726), .ZN(n518) );
  INV_X1 U612 ( .A(KEYINPUT44), .ZN(n527) );
  NAND2_X1 U613 ( .A1(n527), .A2(KEYINPUT90), .ZN(n517) );
  NAND2_X1 U614 ( .A1(n643), .A2(n644), .ZN(n519) );
  XNOR2_X1 U615 ( .A(n520), .B(KEYINPUT33), .ZN(n672) );
  NOR2_X1 U616 ( .A1(n531), .A2(n672), .ZN(n521) );
  XNOR2_X1 U617 ( .A(n521), .B(KEYINPUT34), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n533), .A2(n522), .ZN(n550) );
  XOR2_X1 U619 ( .A(KEYINPUT80), .B(n550), .Z(n523) );
  NAND2_X1 U620 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U621 ( .A(n525), .B(KEYINPUT35), .ZN(n526) );
  NAND2_X1 U622 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U623 ( .A1(n546), .A2(n529), .ZN(n652) );
  NOR2_X1 U624 ( .A1(n652), .A2(n531), .ZN(n530) );
  XNOR2_X1 U625 ( .A(n530), .B(KEYINPUT31), .ZN(n628) );
  NOR2_X1 U626 ( .A1(n531), .A2(n546), .ZN(n532) );
  NAND2_X1 U627 ( .A1(n628), .A2(n609), .ZN(n536) );
  NOR2_X1 U628 ( .A1(n533), .A2(n534), .ZN(n617) );
  INV_X1 U629 ( .A(n617), .ZN(n629) );
  NAND2_X1 U630 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U631 ( .A(n535), .B(KEYINPUT102), .ZN(n626) );
  NAND2_X1 U632 ( .A1(n629), .A2(n626), .ZN(n657) );
  AND2_X1 U633 ( .A1(n536), .A2(n657), .ZN(n540) );
  NOR2_X1 U634 ( .A1(n578), .A2(n537), .ZN(n538) );
  NAND2_X1 U635 ( .A1(n644), .A2(n538), .ZN(n539) );
  XNOR2_X1 U636 ( .A(KEYINPUT103), .B(n539), .ZN(n725) );
  NOR2_X1 U637 ( .A1(n540), .A2(n725), .ZN(n541) );
  NOR2_X1 U638 ( .A1(G900), .A2(n543), .ZN(n544) );
  NOR2_X1 U639 ( .A1(n545), .A2(n544), .ZN(n552) );
  INV_X1 U640 ( .A(n596), .ZN(n548) );
  NOR2_X1 U641 ( .A1(n566), .A2(n548), .ZN(n549) );
  XNOR2_X1 U642 ( .A(n549), .B(KEYINPUT107), .ZN(n551) );
  XNOR2_X1 U643 ( .A(n622), .B(KEYINPUT83), .ZN(n560) );
  NOR2_X1 U644 ( .A1(n644), .A2(n552), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n553), .A2(n643), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n554), .A2(n579), .ZN(n555) );
  XNOR2_X1 U647 ( .A(n555), .B(KEYINPUT28), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n557), .A2(n385), .ZN(n572) );
  NOR2_X1 U649 ( .A1(n558), .A2(n572), .ZN(n623) );
  NAND2_X1 U650 ( .A1(n623), .A2(n657), .ZN(n562) );
  NAND2_X1 U651 ( .A1(KEYINPUT47), .A2(n562), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U653 ( .A(KEYINPUT82), .B(n561), .Z(n565) );
  NOR2_X1 U654 ( .A1(KEYINPUT47), .A2(n562), .ZN(n563) );
  XNOR2_X1 U655 ( .A(n563), .B(KEYINPUT77), .ZN(n564) );
  NAND2_X1 U656 ( .A1(n565), .A2(n564), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n596), .B(KEYINPUT38), .ZN(n658) );
  NOR2_X1 U658 ( .A1(n566), .A2(n658), .ZN(n568) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n568), .B(n567), .ZN(n592) );
  INV_X1 U661 ( .A(n626), .ZN(n624) );
  NAND2_X1 U662 ( .A1(n592), .A2(n624), .ZN(n570) );
  INV_X1 U663 ( .A(KEYINPUT40), .ZN(n569) );
  XNOR2_X1 U664 ( .A(n570), .B(n569), .ZN(n729) );
  INV_X1 U665 ( .A(n729), .ZN(n574) );
  INV_X1 U666 ( .A(n661), .ZN(n571) );
  NAND2_X1 U667 ( .A1(n574), .A2(n727), .ZN(n575) );
  XNOR2_X1 U668 ( .A(n575), .B(KEYINPUT46), .ZN(n576) );
  NOR2_X1 U669 ( .A1(n577), .A2(n576), .ZN(n588) );
  INV_X1 U670 ( .A(n578), .ZN(n580) );
  XNOR2_X1 U671 ( .A(n581), .B(KEYINPUT105), .ZN(n582) );
  NOR2_X1 U672 ( .A1(n626), .A2(n582), .ZN(n583) );
  XNOR2_X1 U673 ( .A(KEYINPUT106), .B(n583), .ZN(n584) );
  INV_X1 U674 ( .A(n584), .ZN(n594) );
  NOR2_X1 U675 ( .A1(n594), .A2(n585), .ZN(n586) );
  XNOR2_X1 U676 ( .A(KEYINPUT36), .B(n586), .ZN(n587) );
  NAND2_X1 U677 ( .A1(n587), .A2(n595), .ZN(n633) );
  NAND2_X1 U678 ( .A1(n588), .A2(n633), .ZN(n591) );
  XOR2_X1 U679 ( .A(KEYINPUT48), .B(KEYINPUT71), .Z(n589) );
  NAND2_X1 U680 ( .A1(n617), .A2(n592), .ZN(n634) );
  INV_X1 U681 ( .A(n593), .ZN(n663) );
  INV_X1 U682 ( .A(n635), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n602), .A2(n598), .ZN(n600) );
  XOR2_X1 U684 ( .A(KEYINPUT62), .B(KEYINPUT91), .Z(n604) );
  NOR2_X1 U685 ( .A1(n626), .A2(n609), .ZN(n607) );
  XNOR2_X1 U686 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U688 ( .A(G104), .B(n608), .ZN(G6) );
  NOR2_X1 U689 ( .A1(n629), .A2(n609), .ZN(n614) );
  XOR2_X1 U690 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n611) );
  XNOR2_X1 U691 ( .A(G107), .B(KEYINPUT26), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT110), .B(n612), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n614), .B(n613), .ZN(G9) );
  XOR2_X1 U695 ( .A(G110), .B(n615), .Z(n616) );
  XNOR2_X1 U696 ( .A(KEYINPUT112), .B(n616), .ZN(G12) );
  XOR2_X1 U697 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n619) );
  NAND2_X1 U698 ( .A1(n623), .A2(n617), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n619), .B(n618), .ZN(n621) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT113), .Z(n620) );
  XNOR2_X1 U701 ( .A(n621), .B(n620), .ZN(G30) );
  XOR2_X1 U702 ( .A(G143), .B(n622), .Z(G45) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n625), .B(G146), .ZN(G48) );
  NOR2_X1 U705 ( .A1(n626), .A2(n628), .ZN(n627) );
  XOR2_X1 U706 ( .A(G113), .B(n627), .Z(G15) );
  NOR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n631) );
  XNOR2_X1 U708 ( .A(G116), .B(KEYINPUT115), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(G18) );
  XOR2_X1 U710 ( .A(G125), .B(KEYINPUT37), .Z(n632) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G134), .B(n634), .ZN(G36) );
  XOR2_X1 U713 ( .A(n635), .B(G140), .Z(G42) );
  XOR2_X1 U714 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n678) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT85), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n719), .A2(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U718 ( .A(KEYINPUT50), .B(n642), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U720 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT116), .B(n647), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n546), .A2(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U726 ( .A(KEYINPUT51), .B(n653), .Z(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U728 ( .A(KEYINPUT118), .B(n656), .Z(n668) );
  INV_X1 U729 ( .A(n657), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n672), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n669), .B(KEYINPUT52), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U740 ( .A(KEYINPUT119), .B(n676), .ZN(n677) );
  XNOR2_X1 U741 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT57), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n682), .B(n681), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n697), .A2(G469), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n699), .A2(n685), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n697), .A2(G475), .ZN(n689) );
  INV_X1 U748 ( .A(KEYINPUT59), .ZN(n686) );
  XNOR2_X1 U749 ( .A(KEYINPUT60), .B(n691), .ZN(G60) );
  NAND2_X1 U750 ( .A1(n697), .A2(G478), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n692), .B(KEYINPUT122), .ZN(n693) );
  XNOR2_X1 U752 ( .A(KEYINPUT124), .B(n700), .ZN(G66) );
  NAND2_X1 U753 ( .A1(n448), .A2(n701), .ZN(n705) );
  NAND2_X1 U754 ( .A1(G953), .A2(G224), .ZN(n702) );
  XNOR2_X1 U755 ( .A(KEYINPUT61), .B(n702), .ZN(n703) );
  NAND2_X1 U756 ( .A1(n703), .A2(G898), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n711) );
  XOR2_X1 U758 ( .A(n706), .B(n707), .Z(n709) );
  NOR2_X1 U759 ( .A1(G898), .A2(n448), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U762 ( .A(KEYINPUT125), .B(n712), .Z(G69) );
  XOR2_X1 U763 ( .A(n714), .B(n713), .Z(n720) );
  XOR2_X1 U764 ( .A(G227), .B(n720), .Z(n715) );
  NAND2_X1 U765 ( .A1(n715), .A2(G900), .ZN(n716) );
  XOR2_X1 U766 ( .A(KEYINPUT126), .B(n716), .Z(n717) );
  NOR2_X1 U767 ( .A1(n448), .A2(n717), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT127), .ZN(n723) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n721), .A2(n448), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n723), .A2(n722), .ZN(G72) );
  XNOR2_X1 U772 ( .A(G122), .B(n724), .ZN(G24) );
  XOR2_X1 U773 ( .A(G101), .B(n725), .Z(G3) );
  XOR2_X1 U774 ( .A(n726), .B(G119), .Z(G21) );
  XOR2_X1 U775 ( .A(G137), .B(n728), .Z(G39) );
  XOR2_X1 U776 ( .A(G131), .B(n729), .Z(G33) );
endmodule

