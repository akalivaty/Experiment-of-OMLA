//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G116), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n187), .A2(new_n190), .ZN(new_n195));
  INV_X1    g009(.A(new_n191), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT66), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(G143), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n210), .A3(new_n205), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G134), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n222), .A3(new_n218), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n201), .A2(new_n203), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n206), .B2(G146), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n225), .A2(new_n206), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n205), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(G146), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n237));
  OAI22_X1  g051(.A1(new_n235), .A2(G143), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n238), .B2(new_n231), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n212), .B(new_n224), .C1(new_n233), .C2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(new_n204), .A3(G128), .A4(new_n207), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n204), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n245), .B2(new_n229), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n217), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n247), .B2(new_n214), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n223), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n199), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n246), .B2(new_n249), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT71), .B1(new_n240), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n240), .A2(KEYINPUT71), .A3(new_n257), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n254), .B(new_n255), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n240), .A2(new_n250), .A3(new_n199), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT26), .B(G101), .Z(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n264), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n268), .B(new_n269), .Z(new_n270));
  NOR2_X1   g084(.A1(new_n259), .A2(new_n258), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT67), .B1(new_n229), .B2(new_n232), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n238), .A2(new_n234), .A3(new_n231), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n272), .A2(new_n273), .B1(new_n209), .B2(new_n211), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n224), .B1(new_n246), .B2(new_n249), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n198), .B1(new_n275), .B2(new_n252), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT72), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n262), .A2(new_n263), .A3(new_n270), .A4(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n277), .A2(new_n270), .A3(new_n261), .A4(new_n260), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n240), .A2(new_n250), .A3(new_n199), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n199), .B1(new_n240), .B2(new_n250), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT28), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n261), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n270), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n278), .A2(new_n280), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT32), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT32), .B1(new_n289), .B2(new_n290), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n261), .A3(new_n260), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n287), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n270), .A3(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT74), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n295), .B2(new_n287), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n297), .A2(new_n298), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT75), .B1(new_n308), .B2(G472), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n303), .B2(new_n304), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT74), .B(new_n299), .C1(new_n287), .C2(new_n295), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT75), .B(G472), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n294), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(KEYINPUT16), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n200), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n316), .B(G146), .C1(KEYINPUT16), .C2(new_n318), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n190), .B2(G128), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n324), .B(new_n325), .C1(G119), .C2(new_n243), .ZN(new_n326));
  XNOR2_X1  g140(.A(G119), .B(G128), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT24), .B(G110), .Z(new_n328));
  AOI22_X1  g142(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n235), .A2(new_n315), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n321), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT76), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n334), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(G234), .B2(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n206), .A2(KEYINPUT80), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT80), .B(G143), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n352), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT18), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n222), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n332), .B1(new_n200), .B2(new_n315), .ZN(new_n360));
  OAI21_X1  g174(.A(G131), .B1(new_n354), .B2(new_n356), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n359), .B(new_n360), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G113), .B(G122), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n222), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT17), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n320), .B(new_n321), .C1(new_n361), .C2(new_n367), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n362), .B(new_n365), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n361), .A2(new_n367), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n320), .A4(new_n321), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n365), .B1(new_n374), .B2(new_n362), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n341), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT82), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n378), .B(new_n341), .C1(new_n372), .C2(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G475), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT19), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n315), .B(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n321), .B1(new_n382), .B2(new_n225), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT81), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n366), .A2(new_n361), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n321), .B(new_n386), .C1(new_n382), .C2(new_n225), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n365), .B1(new_n388), .B2(new_n362), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n372), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT20), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n394), .B(new_n391), .C1(new_n372), .C2(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n380), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT13), .B1(new_n243), .B2(G143), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n217), .ZN(new_n399));
  XNOR2_X1  g213(.A(G128), .B(G143), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n188), .A2(G122), .ZN(new_n402));
  INV_X1    g216(.A(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G116), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT83), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n402), .B2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n401), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n187), .A2(KEYINPUT14), .A3(new_n403), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n406), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n400), .A2(G134), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(G134), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n410), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT9), .B(G234), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n419), .A2(new_n345), .A3(G953), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n410), .B(new_n420), .C1(new_n414), .C2(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G478), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n424), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n397), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  INV_X1    g243(.A(new_n224), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n364), .A2(G107), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n364), .A2(G107), .ZN(new_n433));
  OAI21_X1  g247(.A(G101), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT3), .B1(new_n364), .B2(G107), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT3), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n406), .A3(G104), .ZN(new_n437));
  INV_X1    g251(.A(G101), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .A4(new_n431), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n246), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n242), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n204), .A2(new_n207), .B1(G128), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n430), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n440), .A2(KEYINPUT10), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n246), .A2(new_n449), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n435), .A2(new_n437), .A3(new_n431), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(G101), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(G101), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT4), .A3(new_n439), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n274), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n457), .A3(new_n430), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G140), .ZN(new_n459));
  INV_X1    g273(.A(G227), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n448), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n451), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n224), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(new_n458), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n429), .B(new_n341), .C1(new_n465), .C2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n458), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n462), .B1(new_n448), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n463), .A3(new_n458), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(G469), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n429), .A2(new_n341), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G221), .B1(new_n419), .B2(G902), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n477), .B(KEYINPUT77), .Z(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n266), .A2(G224), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G125), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n274), .A2(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n246), .A2(G125), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n481), .C1(new_n483), .C2(new_n274), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n198), .A2(new_n454), .A3(new_n456), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n189), .A2(new_n191), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n191), .ZN(new_n493));
  INV_X1    g307(.A(G113), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n194), .A3(new_n440), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G110), .B(G122), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n497), .A3(new_n499), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G210), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n484), .A2(new_n486), .B1(new_n508), .B2(new_n482), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n499), .B(KEYINPUT8), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n194), .A2(new_n440), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n189), .A2(KEYINPUT5), .A3(new_n191), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n495), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n440), .B1(new_n496), .B2(new_n194), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n482), .A2(new_n508), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n485), .B(new_n516), .C1(new_n483), .C2(new_n274), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n509), .A2(new_n502), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n506), .A2(new_n341), .A3(new_n507), .A4(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n507), .B(KEYINPUT79), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n341), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n506), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G952), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G953), .ZN(new_n527));
  NAND2_X1  g341(.A1(G234), .A2(G237), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(G902), .A3(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT21), .B(G898), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G214), .B1(G237), .B2(G902), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR4_X1   g351(.A1(new_n428), .A2(new_n480), .A3(new_n525), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n314), .A2(new_n351), .A3(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT84), .B(G101), .Z(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(G3));
  NAND2_X1  g355(.A1(new_n289), .A2(new_n341), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n288), .B1(new_n279), .B2(KEYINPUT31), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n290), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n548));
  OR3_X1    g362(.A1(new_n424), .A2(new_n548), .A3(G478), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n424), .B2(G478), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n422), .A2(new_n423), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT33), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n422), .A2(new_n553), .A3(new_n423), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n425), .A2(G902), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n549), .A2(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n397), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n507), .A4(new_n506), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n519), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n507), .B1(new_n523), .B2(new_n506), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n536), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n559), .A2(new_n534), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n480), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n547), .A2(new_n565), .A3(new_n351), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G104), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G6));
  INV_X1    g384(.A(new_n427), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n397), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n572), .A2(KEYINPUT88), .A3(new_n534), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n380), .A2(new_n396), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n427), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n576), .B2(new_n535), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n573), .A2(new_n577), .A3(new_n564), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n351), .A3(new_n566), .A4(new_n547), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G107), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G9));
  INV_X1    g395(.A(new_n348), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n334), .A2(KEYINPUT89), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n334), .A2(KEYINPUT89), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n585), .A2(KEYINPUT36), .A3(new_n338), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(KEYINPUT36), .B2(new_n338), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n347), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n547), .A2(new_n538), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT37), .B(G110), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G12));
  NAND2_X1  g406(.A1(new_n566), .A2(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT90), .B(G900), .Z(new_n595));
  AOI21_X1  g409(.A(new_n530), .B1(new_n532), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n576), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n564), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n314), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n310), .B2(new_n311), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n312), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n593), .B1(new_n606), .B2(new_n294), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT91), .A3(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT92), .B(G128), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G30));
  XOR2_X1   g425(.A(new_n596), .B(KEYINPUT39), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n566), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT95), .Z(new_n614));
  OR2_X1    g428(.A1(new_n614), .A2(KEYINPUT40), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n287), .B1(new_n281), .B2(new_n282), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT94), .Z(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n279), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n618), .B2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n294), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n614), .A2(KEYINPUT40), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n525), .B(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n536), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n427), .B1(new_n380), .B2(new_n396), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR4_X1   g441(.A1(new_n624), .A2(new_n625), .A3(new_n589), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n615), .A2(new_n620), .A3(new_n621), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G143), .ZN(G45));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n558), .A2(new_n597), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n632), .B2(new_n564), .ZN(new_n633));
  INV_X1    g447(.A(new_n564), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(KEYINPUT96), .A3(new_n558), .A4(new_n597), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n607), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  INV_X1    g452(.A(new_n468), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n448), .B2(new_n464), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n341), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G469), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n479), .A3(new_n469), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n314), .A2(new_n351), .A3(new_n565), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT41), .B(G113), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G15));
  NAND4_X1  g461(.A1(new_n314), .A2(new_n351), .A3(new_n578), .A4(new_n644), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G116), .ZN(G18));
  NAND2_X1  g463(.A1(new_n589), .A2(new_n535), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n650), .A2(new_n643), .A3(new_n428), .A4(new_n564), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n314), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G119), .ZN(G21));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n270), .B1(new_n286), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n283), .A2(KEYINPUT97), .A3(new_n285), .ZN(new_n656));
  AOI22_X1  g470(.A1(KEYINPUT31), .A2(new_n279), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n278), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n280), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n290), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n351), .A3(new_n543), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n642), .A2(new_n479), .A3(new_n469), .A4(new_n535), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT99), .B1(new_n564), .B2(new_n627), .ZN(new_n665));
  INV_X1    g479(.A(new_n507), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n524), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n561), .A3(new_n519), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n625), .B1(new_n520), .B2(KEYINPUT85), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .A4(new_n626), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n664), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n663), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G122), .ZN(G24));
  NAND3_X1  g488(.A1(new_n662), .A2(new_n543), .A3(new_n589), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n662), .A2(KEYINPUT100), .A3(new_n543), .A4(new_n589), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n632), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n644), .A2(new_n634), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n525), .A2(new_n536), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n480), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n480), .A2(new_n688), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n314), .A2(new_n351), .A3(new_n692), .A4(new_n680), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT32), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n546), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n291), .B1(new_n293), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n350), .B1(new_n699), .B2(new_n606), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n690), .A2(new_n632), .A3(new_n691), .A4(new_n685), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n685), .A2(new_n693), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n222), .ZN(G33));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n598), .B(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n314), .A2(new_n351), .A3(new_n692), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n350), .B1(new_n606), .B2(new_n294), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n692), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G134), .ZN(G36));
  NOR2_X1   g526(.A1(new_n575), .A2(new_n557), .ZN(new_n713));
  NOR2_X1   g527(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n714));
  AND2_X1   g528(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n713), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n589), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n547), .ZN(new_n719));
  OR3_X1    g533(.A1(new_n719), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT45), .B1(new_n471), .B2(new_n472), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n429), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n471), .A2(KEYINPUT45), .A3(new_n472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n475), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(KEYINPUT46), .A3(new_n475), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n469), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n479), .A3(new_n612), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT105), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n686), .B1(new_n719), .B2(KEYINPUT44), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT107), .B1(new_n719), .B2(KEYINPUT44), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n720), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n729), .B(new_n479), .C1(KEYINPUT108), .C2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n729), .A2(new_n479), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n680), .A2(new_n350), .A3(new_n687), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n740), .A2(new_n314), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n317), .ZN(G42));
  NOR3_X1   g557(.A1(new_n480), .A2(new_n525), .A3(new_n537), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n559), .A2(new_n572), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n547), .A2(new_n351), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n539), .A2(new_n590), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n692), .A2(new_n680), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n686), .A2(new_n428), .A3(new_n596), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n750), .A2(new_n679), .B1(new_n607), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n711), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n693), .A2(new_n685), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n700), .A2(new_n701), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n314), .A2(new_n651), .B1(new_n663), .B2(new_n672), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(new_n645), .A3(new_n648), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT109), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n645), .A3(new_n648), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n702), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n749), .B1(new_n678), .B2(new_n677), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n607), .A2(new_n751), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n747), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n765), .A3(new_n766), .A4(new_n711), .ZN(new_n767));
  INV_X1    g581(.A(new_n589), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n566), .A3(new_n597), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n665), .B2(new_n671), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n607), .A2(new_n636), .B1(new_n770), .B2(new_n620), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT91), .B1(new_n607), .B2(new_n599), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n695), .A2(new_n291), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n605), .B2(new_n312), .ZN(new_n774));
  INV_X1    g588(.A(new_n599), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n774), .A2(new_n601), .A3(new_n775), .A4(new_n593), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n771), .B(new_n683), .C1(new_n772), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n609), .A2(KEYINPUT52), .A3(new_n683), .A4(new_n771), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n760), .A2(new_n767), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n781), .B2(KEYINPUT110), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n760), .A2(new_n767), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n783), .B(KEYINPUT54), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT111), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n779), .A2(new_n780), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n785), .B1(new_n792), .B2(new_n784), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT112), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n794), .A2(new_n795), .A3(new_n788), .A4(new_n753), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n782), .A2(new_n788), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n789), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n793), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT54), .A4(new_n783), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n530), .A2(new_n717), .A3(new_n644), .A4(new_n687), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n700), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT48), .Z(new_n807));
  INV_X1    g621(.A(new_n620), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n643), .A2(new_n686), .A3(new_n350), .A4(new_n529), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n558), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n663), .A2(new_n530), .A3(new_n717), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n810), .B(new_n527), .C1(new_n681), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n644), .A2(new_n625), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n623), .B1(KEYINPUT114), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n642), .A2(new_n469), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n478), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n740), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n687), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n811), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n397), .A2(new_n808), .A3(new_n557), .A4(new_n809), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n679), .B2(new_n805), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n819), .B1(new_n818), .B2(new_n811), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n813), .B1(new_n830), .B2(KEYINPUT51), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n832), .B(KEYINPUT51), .C1(new_n811), .C2(new_n824), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n791), .A2(new_n800), .A3(new_n804), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n526), .A2(new_n266), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n821), .B(KEYINPUT49), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n351), .A2(new_n479), .A3(new_n536), .A4(new_n713), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n808), .A2(new_n624), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(G75));
  NOR2_X1   g661(.A1(new_n266), .A2(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n797), .A2(new_n799), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(G902), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n852), .B2(G210), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n503), .A2(new_n505), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(new_n489), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT55), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n849), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT56), .B1(new_n857), .B2(KEYINPUT118), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(KEYINPUT118), .B2(new_n857), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n521), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  INV_X1    g676(.A(new_n521), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n860), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n858), .A2(new_n865), .ZN(G51));
  NOR2_X1   g680(.A1(new_n851), .A2(new_n724), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n474), .B(KEYINPUT119), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT57), .Z(new_n869));
  AND3_X1   g683(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n640), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT120), .B1(new_n873), .B2(new_n848), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n875));
  INV_X1    g689(.A(new_n640), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n800), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n878), .B2(new_n869), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n875), .B(new_n849), .C1(new_n879), .C2(new_n867), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n852), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(new_n390), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n390), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n848), .ZN(G60));
  XNOR2_X1  g699(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n425), .A2(new_n341), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n886), .B(new_n887), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n804), .A2(new_n800), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n801), .A2(new_n793), .B1(KEYINPUT53), .B2(new_n782), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n803), .B1(new_n891), .B2(KEYINPUT54), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n555), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n888), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n848), .B1(new_n878), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(KEYINPUT122), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n791), .A2(new_n800), .A3(new_n804), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n555), .B1(new_n900), .B2(new_n889), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n896), .B1(new_n870), .B2(new_n871), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n849), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n898), .A2(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n797), .B2(new_n799), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n340), .B(KEYINPUT123), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n588), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n848), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n908), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n913), .B(new_n916), .ZN(G66));
  INV_X1    g731(.A(new_n533), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n266), .B1(new_n918), .B2(G224), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n761), .A2(new_n747), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(new_n266), .ZN(new_n922));
  INV_X1    g736(.A(G898), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n854), .B1(new_n923), .B2(G953), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n922), .B(new_n924), .ZN(G69));
  INV_X1    g739(.A(new_n614), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n926), .A2(new_n709), .A3(new_n687), .A4(new_n745), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n734), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n734), .A2(KEYINPUT125), .A3(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n742), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n629), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n609), .A2(new_n637), .A3(new_n683), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n933), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n932), .A2(new_n266), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n259), .A2(new_n258), .B1(new_n275), .B2(new_n252), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(new_n382), .Z(new_n939));
  NAND3_X1  g753(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n939), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n460), .A2(G900), .A3(G953), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n665), .A2(new_n671), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n731), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n742), .B1(new_n945), .B2(new_n700), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n756), .A3(new_n711), .ZN(new_n947));
  INV_X1    g761(.A(new_n734), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n948), .A2(new_n949), .A3(new_n934), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n948), .B2(new_n934), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n942), .B(new_n943), .C1(new_n952), .C2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n941), .A2(new_n953), .ZN(G72));
  NOR2_X1   g768(.A1(new_n295), .A2(new_n270), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n920), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n932), .A2(new_n920), .A3(new_n935), .A4(new_n936), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n958), .ZN(new_n962));
  INV_X1    g776(.A(new_n295), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n287), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n848), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n959), .A3(new_n955), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n891), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n960), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G57));
endmodule


