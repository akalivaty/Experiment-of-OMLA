//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1190, new_n1191,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  MUX2_X1   g039(.A(new_n463), .B(new_n464), .S(G2105), .Z(G160));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n462), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT69), .Z(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n468), .A2(new_n470), .A3(G126), .ZN(new_n484));
  NAND2_X1  g059(.A1(G114), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n472), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G102), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n483), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n485), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(G126), .ZN(new_n492));
  OAI211_X1 g067(.A(KEYINPUT70), .B(new_n488), .C1(new_n492), .C2(new_n472), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n472), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(G75), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(G651), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(G651), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(new_n506), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G88), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT73), .B(G651), .C1(new_n507), .C2(new_n508), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n511), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND4_X1  g101(.A1(new_n517), .A2(new_n520), .A3(G89), .A4(new_n518), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n517), .A2(G51), .A3(G543), .A4(new_n518), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n515), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n519), .A2(G90), .A3(new_n520), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n522), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G81), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n519), .A2(new_n520), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n522), .A2(G43), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n504), .B2(new_n506), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND4_X1  g128(.A1(new_n517), .A2(new_n520), .A3(G91), .A4(new_n518), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n517), .A2(G53), .A3(G543), .A4(new_n518), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n515), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(G299));
  XNOR2_X1  g136(.A(new_n532), .B(KEYINPUT76), .ZN(G286));
  NAND3_X1  g137(.A1(new_n519), .A2(G87), .A3(new_n520), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n522), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n504), .B2(new_n506), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n517), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n517), .A2(new_n520), .A3(G86), .A4(new_n518), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n515), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n519), .A2(G85), .A3(new_n520), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(G47), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n517), .A2(new_n520), .A3(G92), .A4(new_n518), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n522), .A2(G54), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n504), .B2(new_n506), .ZN(new_n587));
  AND2_X1   g162(.A1(G79), .A2(G543), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n587), .A2(KEYINPUT78), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(G651), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n584), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n581), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n581), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  XNOR2_X1  g170(.A(G299), .B(KEYINPUT79), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g179(.A1(new_n475), .A2(G123), .B1(G135), .B2(new_n478), .ZN(new_n605));
  NOR2_X1   g180(.A1(G99), .A2(G2105), .ZN(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G2096), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n462), .A2(new_n487), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT13), .B(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(G2443), .B(G2446), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2435), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2438), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n618), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n632), .A2(new_n617), .A3(new_n628), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n633), .A3(G14), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n637), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n641), .B2(new_n638), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(KEYINPUT83), .C1(new_n641), .C2(new_n638), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n643), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n637), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n639), .A3(new_n640), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  AND3_X1   g229(.A1(new_n651), .A2(new_n609), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n609), .B1(new_n651), .B2(new_n654), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n636), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n649), .A2(new_n650), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n654), .A3(new_n642), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G2096), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n651), .A2(new_n609), .A3(new_n654), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(G2100), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(new_n684), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G25), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n475), .A2(G119), .B1(G131), .B2(new_n478), .ZN(new_n690));
  OR2_X1    g265(.A1(G95), .A2(G2105), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n691), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n689), .B1(new_n693), .B2(G29), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT35), .B(G1991), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G24), .ZN(new_n699));
  INV_X1    g274(.A(G290), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(G1986), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n697), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n698), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n698), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT86), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n710), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n710), .A2(KEYINPUT34), .A3(new_n715), .A4(new_n719), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n706), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT88), .B1(new_n724), .B2(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n722), .A2(new_n723), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(new_n705), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT87), .B1(new_n731), .B2(KEYINPUT36), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n724), .A2(new_n733), .A3(new_n725), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n728), .A2(new_n729), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n688), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n688), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT29), .B(G2090), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n688), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n487), .A2(G103), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n478), .A2(G139), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n472), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n740), .B1(new_n751), .B2(new_n688), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2072), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n698), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n592), .B2(new_n698), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1348), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n698), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n547), .B2(new_n698), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1341), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n688), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n475), .A2(G128), .B1(G140), .B2(new_n478), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n762), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n756), .A2(new_n759), .A3(new_n769), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT90), .Z(new_n771));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI22_X1  g351(.A1(G160), .A2(G29), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n772), .B2(new_n776), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2084), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT31), .B(G11), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT95), .B(G28), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT30), .Z(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(G29), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT26), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n475), .B2(G129), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n487), .A2(G105), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n478), .A2(G141), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G32), .B(new_n789), .S(G29), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT27), .B(G1996), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n608), .A2(new_n688), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n783), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n752), .A2(G2072), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n688), .A2(G27), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n688), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n698), .A2(G20), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G299), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n698), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1956), .ZN(new_n805));
  NAND2_X1  g380(.A1(G171), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G5), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G1966), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n532), .A2(G16), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G21), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n809), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n807), .A2(new_n808), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n805), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n794), .A2(new_n795), .A3(new_n799), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n771), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n735), .A2(new_n739), .A3(new_n753), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n813), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(G1966), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(G311));
  OR2_X1    g397(.A1(new_n771), .A2(new_n817), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n732), .A2(new_n734), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n726), .B(new_n727), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n821), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n739), .A4(new_n753), .ZN(G150));
  AND2_X1   g403(.A1(new_n520), .A2(G67), .ZN(new_n829));
  AND2_X1   g404(.A1(G80), .A2(G543), .ZN(new_n830));
  OAI21_X1  g405(.A(G651), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n522), .A2(G55), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT97), .B(G93), .Z(new_n833));
  NAND3_X1  g408(.A1(new_n519), .A2(new_n520), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n547), .A2(new_n835), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(new_n831), .A3(new_n832), .A4(new_n834), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n592), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n837), .B1(new_n845), .B2(G860), .ZN(G145));
  XNOR2_X1  g421(.A(new_n608), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n475), .A2(G130), .B1(G142), .B2(new_n478), .ZN(new_n849));
  NOR2_X1   g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n693), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n613), .Z(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(KEYINPUT99), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n488), .B1(new_n492), .B2(new_n472), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n496), .A2(new_n497), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n766), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n789), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n751), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n859), .A2(new_n789), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n789), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n750), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n848), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n861), .B(new_n864), .C1(new_n854), .C2(KEYINPUT99), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n854), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n853), .B(new_n613), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT98), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n870), .A2(new_n872), .A3(new_n864), .A4(new_n861), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n869), .A3(new_n854), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(new_n848), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT100), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(KEYINPUT40), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(G395));
  INV_X1    g459(.A(G868), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n601), .B(new_n841), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n584), .A2(new_n585), .A3(new_n591), .ZN(new_n887));
  NAND2_X1  g462(.A1(G299), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(G299), .A2(new_n887), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n803), .A2(new_n592), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n888), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n886), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n712), .A2(G305), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n712), .A2(G305), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n700), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n712), .A2(G305), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(G290), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G303), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(new_n909), .A3(G166), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n903), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n900), .A2(new_n915), .A3(new_n902), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n885), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n835), .A2(new_n885), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n917), .A2(KEYINPUT101), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n921));
  INV_X1    g496(.A(new_n916), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n915), .B1(new_n900), .B2(new_n902), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n924), .B2(new_n918), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n920), .A2(new_n925), .ZN(G295));
  NOR3_X1   g501(.A1(new_n917), .A2(KEYINPUT102), .A3(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n924), .B2(new_n918), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n835), .B(new_n839), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT76), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n532), .B(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(G301), .ZN(new_n935));
  NAND2_X1  g510(.A1(G301), .A2(G168), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n932), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G286), .A2(G171), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n841), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n895), .A4(new_n897), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n895), .A2(new_n938), .A3(new_n897), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT103), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n891), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n945), .A3(new_n915), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n944), .A2(KEYINPUT103), .B1(new_n891), .B2(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n915), .B1(new_n951), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n931), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n947), .A2(new_n944), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n913), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n949), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n931), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n950), .B2(new_n952), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n948), .A2(new_n955), .A3(new_n931), .A4(new_n949), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(KEYINPUT104), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n960), .A2(KEYINPUT104), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n963), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g539(.A(new_n766), .B(G2067), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n856), .B2(new_n857), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G160), .A2(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT105), .B1(new_n965), .B2(new_n970), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n789), .B(G1996), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n970), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n693), .B(new_n696), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(G290), .B(G1986), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n970), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(G299), .B(KEYINPUT57), .Z(new_n983));
  OAI211_X1 g558(.A(KEYINPUT45), .B(new_n966), .C1(new_n856), .C2(new_n857), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n484), .A2(new_n485), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G2105), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(new_n496), .A3(new_n497), .A4(new_n488), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n988), .A2(new_n989), .A3(KEYINPUT45), .A4(new_n966), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n969), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n499), .A2(new_n966), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT56), .B(G2072), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(KEYINPUT115), .A3(new_n994), .A4(new_n995), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1956), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n966), .C1(new_n856), .C2(new_n857), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n988), .B2(new_n966), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n969), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1001), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n983), .B1(new_n1000), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n998), .A2(new_n1010), .A3(new_n983), .A4(new_n999), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n969), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1348), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1008), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G2067), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n887), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1011), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n985), .A2(new_n990), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT116), .B(G1996), .Z(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n994), .A3(new_n1008), .A4(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT58), .B(G1341), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(KEYINPUT117), .A3(new_n547), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT59), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(KEYINPUT117), .A3(new_n1029), .A4(new_n547), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n887), .A2(KEYINPUT60), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1028), .A2(new_n1030), .B1(new_n1018), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n1033));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1033), .A2(new_n1034), .B1(KEYINPUT120), .B2(KEYINPUT61), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1012), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1015), .A2(new_n1017), .A3(new_n592), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT60), .B1(new_n1019), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1012), .A2(new_n1039), .A3(KEYINPUT61), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(new_n1036), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1012), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1034), .B1(new_n1042), .B2(new_n1033), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1020), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(G166), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1013), .A2(new_n1014), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1971), .B1(new_n991), .B2(new_n994), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1052), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT109), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1021), .A2(new_n994), .A3(new_n1008), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n709), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1013), .A2(new_n1014), .A3(new_n1053), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(G8), .A4(new_n1052), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G305), .A2(G1981), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT110), .B(G1981), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1016), .A2(new_n1070), .A3(G8), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G288), .A2(new_n1073), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1016), .A2(new_n1074), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n967), .A2(KEYINPUT107), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n969), .B1(new_n1078), .B2(new_n1003), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1079), .A2(new_n1049), .A3(new_n1075), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1072), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1016), .A2(G8), .A3(new_n1076), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT112), .A3(new_n1072), .A4(new_n1077), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1007), .A2(new_n1009), .A3(G2090), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1089), .B2(new_n1055), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1052), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1064), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n1094));
  OR3_X1    g669(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n969), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT122), .B1(new_n1094), .B2(new_n969), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT53), .B1(new_n1097), .B2(G2078), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1097), .B2(G2078), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1095), .A2(new_n1021), .A3(new_n1096), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n808), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1058), .B2(G2078), .ZN(new_n1104));
  XOR2_X1   g679(.A(G301), .B(KEYINPUT54), .Z(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1078), .A2(new_n993), .A3(new_n1003), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1008), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n810), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT113), .B(G2084), .Z(new_n1111));
  NAND3_X1  g686(.A1(new_n1013), .A2(new_n1014), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(G168), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT51), .ZN(new_n1115));
  AOI21_X1  g690(.A(G168), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  OAI211_X1 g692(.A(G8), .B(new_n1113), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(new_n1104), .A3(new_n1102), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1105), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1115), .A2(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1093), .A2(KEYINPUT124), .A3(new_n1106), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1064), .A2(new_n1088), .A3(new_n1092), .A4(new_n1106), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1044), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1072), .A2(new_n1073), .A3(new_n712), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1067), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(G8), .A3(new_n1016), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1082), .B(KEYINPUT111), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n1064), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1061), .A2(G8), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT114), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1061), .A2(new_n1139), .A3(G8), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1091), .A3(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1049), .B(G286), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT111), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1082), .B(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1136), .B1(KEYINPUT63), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1121), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1117), .B1(new_n1113), .B2(G8), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n532), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT51), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1113), .A2(G8), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1150), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(G301), .B1(new_n1127), .B2(KEYINPUT62), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1093), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1146), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n982), .B1(new_n1131), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n980), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n978), .A2(G1996), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT46), .Z(new_n1167));
  OAI21_X1  g742(.A(new_n970), .B1(new_n965), .B2(new_n789), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT47), .Z(new_n1170));
  NOR2_X1   g745(.A1(new_n693), .A2(new_n695), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n977), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n766), .A2(G2067), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(KEYINPUT125), .A3(new_n1174), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n970), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT126), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1177), .A2(new_n1181), .A3(new_n970), .A4(new_n1178), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1165), .B(new_n1170), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1162), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g759(.A(new_n460), .B1(new_n685), .B2(new_n686), .ZN(new_n1186));
  NAND4_X1  g760(.A1(new_n657), .A2(new_n662), .A3(new_n634), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n868), .B2(new_n875), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n1188), .A3(new_n962), .ZN(G225));
  NAND2_X1  g763(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1190));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1191));
  NAND4_X1  g765(.A1(new_n961), .A2(new_n1188), .A3(new_n1191), .A4(new_n962), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1192), .ZN(G308));
endmodule


