//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n202), .A2(new_n203), .B1(new_n204), .B2(KEYINPUT70), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(KEYINPUT70), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n207), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT71), .B1(new_n207), .B2(G120gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G113gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n209), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n204), .A2(new_n203), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n205), .A2(new_n206), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G183gat), .B(G190gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n219), .C1(new_n220), .C2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n218), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n219), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT64), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G169gat), .ZN(new_n229));
  INV_X1    g028(.A(G176gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT23), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n221), .B(new_n228), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT25), .B1(new_n226), .B2(new_n227), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n238), .ZN(new_n244));
  INV_X1    g043(.A(new_n233), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n235), .A2(KEYINPUT26), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n222), .B2(new_n224), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(new_n235), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT27), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G183gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(new_n224), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT68), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(KEYINPUT68), .A3(new_n260), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n256), .A2(new_n258), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n256), .A2(new_n258), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT28), .A4(new_n224), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n255), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n216), .B1(new_n248), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n228), .A2(new_n221), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n240), .B1(new_n244), .B2(new_n245), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n242), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n247), .A2(new_n243), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n216), .ZN(new_n277));
  INV_X1    g076(.A(new_n263), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n269), .B1(new_n278), .B2(new_n261), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n254), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286));
  INV_X1    g085(.A(new_n284), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n282), .B2(KEYINPUT74), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n286), .B(new_n283), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n248), .A2(new_n270), .A3(new_n216), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n277), .B1(new_n276), .B2(new_n280), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n284), .A3(new_n290), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT75), .B1(new_n295), .B2(KEYINPUT34), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n285), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(KEYINPUT76), .B(new_n285), .C1(new_n291), .C2(new_n296), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n271), .A2(new_n281), .A3(new_n287), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT33), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G226gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n274), .A2(new_n275), .B1(new_n279), .B2(new_n254), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n248), .B2(new_n270), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT81), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323));
  INV_X1    g122(.A(G211gat), .ZN(new_n324));
  INV_X1    g123(.A(G218gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT78), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G218gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n332), .B(new_n323), .C1(new_n329), .C2(new_n330), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(KEYINPUT79), .A3(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT80), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n248), .B2(new_n270), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n347), .B2(new_n318), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n322), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n320), .A2(new_n321), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n314), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n348), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n320), .A2(new_n321), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n343), .B(new_n354), .C1(new_n355), .C2(KEYINPUT81), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n351), .A3(new_n313), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n357), .A3(KEYINPUT30), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n349), .A2(new_n352), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n360), .A3(new_n313), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G141gat), .B(G148gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(G155gat), .B2(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G148gat), .ZN(new_n371));
  INV_X1    g170(.A(G148gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G141gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G155gat), .B(G162gat), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n205), .A2(new_n206), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n214), .A2(new_n215), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n389), .B(KEYINPUT83), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n369), .A2(new_n379), .A3(KEYINPUT82), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT3), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n277), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT84), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n388), .A2(new_n391), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n391), .A3(new_n386), .A4(new_n387), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n393), .A2(new_n394), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n277), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n384), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n390), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416));
  INV_X1    g215(.A(new_n414), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n405), .A2(new_n417), .A3(new_n409), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n417), .A4(new_n409), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n362), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G228gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(new_n316), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n346), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n340), .A2(new_n342), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n334), .B2(new_n336), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n380), .B1(new_n427), .B2(KEYINPUT3), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n396), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n406), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(new_n424), .A3(new_n426), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n431), .A2(new_n426), .A3(KEYINPUT86), .A4(new_n424), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G22gat), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G50gat), .ZN(new_n442));
  XOR2_X1   g241(.A(G78gat), .B(G106gat), .Z(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND4_X1  g243(.A1(new_n438), .A2(new_n439), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n439), .B1(new_n436), .B2(new_n437), .ZN(new_n446));
  INV_X1    g245(.A(new_n444), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n436), .A2(new_n437), .ZN(new_n448));
  AOI211_X1 g247(.A(G22gat), .B(new_n429), .C1(new_n434), .C2(new_n435), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n446), .A2(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n309), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n299), .A2(KEYINPUT73), .A3(new_n452), .A4(new_n300), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n310), .A2(new_n422), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  AOI221_X4 g254(.A(KEYINPUT35), .B1(new_n419), .B2(new_n420), .C1(new_n358), .C2(new_n361), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n286), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n295), .A2(KEYINPUT75), .A3(KEYINPUT34), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT76), .B1(new_n460), .B2(new_n285), .ZN(new_n461));
  INV_X1    g260(.A(new_n300), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n309), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n299), .A2(new_n452), .A3(new_n300), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n456), .A2(new_n463), .A3(new_n451), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n299), .A2(new_n452), .A3(new_n300), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n452), .B1(new_n299), .B2(new_n300), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(KEYINPUT91), .A3(new_n451), .A4(new_n456), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n455), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n313), .B1(new_n359), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n350), .B2(new_n343), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n354), .B1(new_n355), .B2(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n343), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT90), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n476), .C1(new_n477), .C2(new_n343), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n474), .A2(new_n475), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n356), .A2(new_n351), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n314), .B1(new_n483), .B2(KEYINPUT37), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n359), .A2(new_n473), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n421), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(new_n486), .A3(new_n487), .A4(new_n357), .ZN(new_n488));
  INV_X1    g287(.A(new_n362), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n391), .B1(new_n388), .B2(new_n398), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT39), .B1(new_n408), .B2(new_n390), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n417), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(KEYINPUT40), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT89), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT40), .B1(new_n492), .B2(new_n494), .ZN(new_n497));
  INV_X1    g296(.A(new_n418), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n488), .A2(new_n500), .A3(new_n451), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n310), .A2(new_n453), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n422), .A2(new_n451), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n463), .A2(new_n507), .A3(new_n464), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n502), .B1(new_n509), .B2(KEYINPUT88), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n310), .B2(new_n453), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT36), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(new_n512), .A3(new_n505), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n472), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT8), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  INV_X1    g321(.A(G92gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n518), .A2(new_n521), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G99gat), .B(G106gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g328(.A1(KEYINPUT8), .A2(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n527), .A3(new_n521), .A4(new_n525), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(KEYINPUT100), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n526), .A2(new_n533), .A3(new_n528), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT98), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  OAI221_X1 g343(.A(new_n537), .B1(new_n541), .B2(new_n542), .C1(new_n538), .C2(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n544), .A2(new_n545), .B1(new_n529), .B2(new_n531), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n535), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n547), .B1(new_n550), .B2(KEYINPUT10), .ZN(new_n551));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT103), .ZN(new_n554));
  INV_X1    g353(.A(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT103), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n551), .A2(new_n560), .A3(new_n552), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n554), .A2(new_n556), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n559), .ZN(new_n563));
  INV_X1    g362(.A(new_n553), .ZN(new_n564));
  INV_X1    g363(.A(new_n556), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT14), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  INV_X1    g375(.A(G43gat), .ZN(new_n577));
  INV_X1    g376(.A(G50gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G43gat), .A2(G50gat), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT93), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n575), .A2(new_n581), .A3(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n575), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n580), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n579), .A2(new_n576), .A3(new_n580), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n585), .A2(KEYINPUT95), .A3(KEYINPUT17), .A4(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n575), .A2(new_n581), .A3(KEYINPUT93), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n590), .B(KEYINPUT17), .C1(new_n592), .C2(new_n582), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n585), .A2(new_n590), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n535), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT101), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n597), .A2(new_n535), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  XOR2_X1   g406(.A(G134gat), .B(G162gat), .Z(new_n608));
  NOR2_X1   g407(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n611), .B(new_n613), .C1(new_n606), .C2(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G8gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G15gat), .B(G22gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT16), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(G1gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n622), .B2(KEYINPUT94), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(G1gat), .B2(new_n620), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI221_X1 g424(.A(new_n622), .B1(KEYINPUT94), .B2(new_n619), .C1(G1gat), .C2(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(KEYINPUT21), .B2(new_n546), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n618), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n629), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n568), .A2(new_n615), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT104), .Z(new_n638));
  AOI21_X1  g437(.A(new_n627), .B1(new_n597), .B2(new_n598), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n596), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n597), .A2(new_n627), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n639), .A2(new_n596), .B1(new_n627), .B2(new_n597), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(KEYINPUT18), .A3(new_n641), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n597), .B(new_n627), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n641), .B(KEYINPUT13), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G169gat), .B(G197gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT12), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(KEYINPUT96), .A3(new_n657), .ZN(new_n661));
  INV_X1    g460(.A(new_n657), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n645), .A2(new_n647), .A3(new_n650), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT97), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n643), .A2(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n647), .A4(new_n662), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n660), .A2(new_n661), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n638), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n516), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n487), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n619), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n489), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n455), .A2(new_n471), .A3(new_n467), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n501), .B1(new_n513), .B2(new_n514), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n489), .A3(new_n669), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G8gat), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n674), .B(new_n679), .C1(new_n686), .C2(new_n678), .ZN(new_n687));
  INV_X1    g486(.A(new_n679), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n678), .B1(new_n677), .B2(new_n685), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT106), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n671), .ZN(new_n692));
  INV_X1    g491(.A(new_n470), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n692), .A2(G15gat), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n504), .A2(new_n508), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1326gat));
  INV_X1    g497(.A(new_n451), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n671), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n668), .A2(new_n636), .A3(new_n567), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n516), .B2(new_n615), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n504), .A2(new_n508), .A3(new_n506), .A4(new_n501), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n680), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n615), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n710));
  OR2_X1    g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n704), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n569), .B1(new_n712), .B2(new_n487), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n421), .A2(G29gat), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n683), .A2(new_n708), .A3(new_n703), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT110), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n683), .B2(new_n708), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n709), .A2(new_n710), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n703), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n421), .ZN(new_n723));
  INV_X1    g522(.A(new_n716), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n715), .B(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n718), .A2(new_n727), .ZN(G1328gat));
  NAND3_X1  g527(.A1(new_n683), .A2(new_n708), .A3(new_n703), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(G36gat), .A3(new_n362), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n722), .B2(new_n362), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(new_n696), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n703), .C1(new_n720), .C2(new_n721), .ZN(new_n735));
  INV_X1    g534(.A(new_n729), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n693), .A2(G43gat), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n735), .A2(G43gat), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n577), .B1(new_n712), .B2(new_n695), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n738), .A2(KEYINPUT47), .B1(new_n739), .B2(new_n741), .ZN(G1330gat));
  NOR2_X1   g541(.A1(new_n451), .A2(new_n578), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n703), .B(new_n743), .C1(new_n720), .C2(new_n721), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n578), .B1(new_n729), .B2(new_n451), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n665), .A2(new_n667), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT96), .B1(new_n651), .B2(new_n657), .ZN(new_n749));
  AOI211_X1 g548(.A(new_n659), .B(new_n662), .C1(new_n666), .C2(new_n647), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n636), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n708), .A4(new_n568), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n707), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n487), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n754), .A2(new_n362), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  NOR3_X1   g561(.A1(new_n754), .A2(G71gat), .A3(new_n693), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n755), .A2(new_n734), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(G71gat), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g565(.A1(new_n754), .A2(new_n451), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT112), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT111), .B(G78gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n421), .A2(G85gat), .A3(new_n568), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n615), .B1(new_n680), .B2(new_n706), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n751), .A2(new_n636), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n773), .B2(new_n774), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n773), .A2(KEYINPUT113), .A3(KEYINPUT51), .A4(new_n774), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(KEYINPUT114), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n771), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n774), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n568), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n720), .B2(new_n721), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n421), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(G1336gat));
  INV_X1    g588(.A(new_n786), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n705), .B2(new_n711), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n523), .B1(new_n791), .B2(new_n489), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n362), .A2(G92gat), .A3(new_n568), .ZN(new_n793));
  AND4_X1   g592(.A1(KEYINPUT51), .A2(new_n707), .A3(new_n708), .A4(new_n774), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n778), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(new_n793), .C1(new_n794), .C2(new_n778), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G92gat), .B1(new_n787), .B2(new_n362), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n781), .B2(new_n793), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1337gat));
  NOR3_X1   g603(.A1(new_n693), .A2(G99gat), .A3(new_n568), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n782), .B2(new_n783), .ZN(new_n806));
  OAI21_X1  g605(.A(G99gat), .B1(new_n787), .B2(new_n696), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1338gat));
  OAI211_X1 g607(.A(new_n699), .B(new_n786), .C1(new_n720), .C2(new_n721), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT116), .B(G106gat), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n451), .A2(G106gat), .A3(new_n568), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n781), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n794), .A2(new_n778), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n809), .A2(new_n810), .B1(new_n816), .B2(new_n812), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n811), .A2(new_n815), .B1(new_n817), .B2(new_n814), .ZN(G1339gat));
  NOR2_X1   g617(.A1(new_n751), .A2(new_n637), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n555), .B(new_n547), .C1(new_n550), .C2(KEYINPUT10), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT10), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n546), .B1(new_n534), .B2(new_n532), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n825), .B2(new_n548), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(KEYINPUT117), .A3(new_n555), .A4(new_n547), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(new_n554), .A3(KEYINPUT54), .A4(new_n561), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n559), .B1(new_n564), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n562), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n829), .B2(new_n831), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n829), .C2(new_n831), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n646), .A2(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n656), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n748), .A2(new_n708), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n748), .A2(new_n567), .A3(new_n841), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n839), .B2(new_n668), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n845), .B2(new_n615), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n820), .B1(new_n846), .B2(new_n636), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n699), .A3(new_n693), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n489), .A2(new_n421), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n207), .A3(new_n668), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n503), .A2(new_n699), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n848), .A2(new_n421), .A3(new_n489), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n751), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n852), .A2(new_n856), .ZN(G1340gat));
  OAI21_X1  g656(.A(G120gat), .B1(new_n851), .B2(new_n568), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT119), .Z(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n211), .A3(new_n567), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n851), .B2(new_n752), .ZN(new_n862));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n863), .A3(new_n636), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1342gat));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n421), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n489), .A2(G134gat), .A3(new_n615), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n853), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n851), .B2(new_n615), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n734), .A2(new_n451), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(new_n362), .A3(new_n866), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n668), .A2(G141gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n695), .A2(new_n421), .A3(new_n489), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n829), .A2(new_n831), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n562), .A3(new_n832), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n844), .B1(new_n668), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n838), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n833), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n842), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n885), .A2(new_n615), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n880), .B1(new_n890), .B2(new_n636), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n751), .A2(new_n834), .A3(new_n883), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n708), .B1(new_n892), .B2(new_n844), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT121), .B(new_n752), .C1(new_n893), .C2(new_n843), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n891), .A2(new_n894), .A3(new_n820), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n451), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n847), .B2(new_n699), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G141gat), .B1(new_n900), .B2(new_n668), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n877), .A2(new_n878), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n847), .A2(new_n699), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n904), .A2(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n905));
  INV_X1    g704(.A(new_n879), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT122), .B(new_n879), .C1(new_n898), .C2(new_n899), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n751), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n875), .A2(new_n876), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n902), .B1(new_n910), .B2(new_n878), .ZN(G1344gat));
  AND2_X1   g710(.A1(new_n847), .A2(new_n897), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n890), .A2(new_n636), .B1(new_n751), .B2(new_n638), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n699), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n567), .B(new_n879), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G148gat), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT59), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n907), .A2(new_n908), .A3(new_n567), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n372), .A2(KEYINPUT59), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n875), .A2(new_n372), .A3(new_n567), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1345gat));
  NAND3_X1  g726(.A1(new_n875), .A2(new_n376), .A3(new_n636), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n907), .A2(new_n636), .A3(new_n908), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n376), .B2(new_n929), .ZN(G1346gat));
  NOR3_X1   g729(.A1(new_n489), .A2(G162gat), .A3(new_n615), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n874), .A2(new_n866), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n907), .A2(new_n708), .A3(new_n908), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n377), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n362), .A2(new_n487), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n849), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n229), .A3(new_n668), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n848), .A2(new_n487), .A3(new_n362), .A4(new_n854), .ZN(new_n938));
  AOI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n751), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1348gat));
  OAI21_X1  g739(.A(G176gat), .B1(new_n936), .B2(new_n568), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n230), .A3(new_n567), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  NOR2_X1   g742(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n944));
  OAI21_X1  g743(.A(G183gat), .B1(new_n936), .B2(new_n752), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n938), .A2(new_n266), .A3(new_n268), .A4(new_n636), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n947), .B(new_n948), .Z(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n936), .B2(new_n615), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n224), .A3(new_n708), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n696), .A2(new_n935), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n912), .A2(new_n914), .ZN(new_n955));
  INV_X1    g754(.A(G197gat), .ZN(new_n956));
  NOR4_X1   g755(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n668), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n696), .A2(new_n958), .A3(new_n489), .A4(new_n699), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(new_n421), .A3(new_n847), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n696), .A2(new_n489), .A3(new_n699), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n751), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n957), .B1(new_n965), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n568), .A2(G204gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n567), .B1(new_n912), .B2(new_n914), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n954), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n968), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT62), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(G1353gat));
  NOR2_X1   g773(.A1(new_n954), .A2(new_n955), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n324), .B1(new_n975), .B2(new_n636), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT63), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n752), .A2(G211gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n962), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(new_n615), .B1(new_n326), .B2(new_n328), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n975), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n964), .A2(new_n708), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(new_n325), .ZN(G1355gat));
endmodule


