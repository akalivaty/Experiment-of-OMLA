//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n435, new_n441, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(new_n435));
  INV_X1    g010(.A(new_n435), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g028(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n466), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n472), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n463), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n465), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(G2104), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n481), .B(new_n484), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT71), .B1(new_n465), .B2(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n465), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n502), .A3(G138), .A4(new_n465), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT72), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n522), .A2(new_n524), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT7), .Z(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n528), .B1(new_n531), .B2(new_n510), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n509), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n509), .A2(new_n518), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(G52), .B2(new_n525), .ZN(G171));
  NAND2_X1  g118(.A1(new_n539), .A2(G81), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n512), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n505), .B1(new_n518), .B2(new_n521), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n547), .A2(G43), .A3(new_n524), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT74), .Z(G188));
  NAND3_X1  g132(.A1(new_n522), .A2(new_n524), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n547), .A2(new_n561), .A3(G53), .A4(new_n524), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n509), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n539), .A2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n563), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  AND3_X1   g147(.A1(new_n526), .A2(KEYINPUT75), .A3(new_n532), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n526), .B2(new_n532), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n525), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n539), .A2(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n509), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(G651), .B1(new_n523), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n539), .A2(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  INV_X1    g164(.A(G72), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n509), .A2(new_n589), .B1(new_n590), .B2(new_n505), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI221_X1 g168(.A(KEYINPUT76), .B1(new_n590), .B2(new_n505), .C1(new_n509), .C2(new_n589), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G651), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n593), .A2(new_n597), .A3(new_n594), .A4(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n539), .A2(G85), .ZN(new_n599));
  INV_X1    g174(.A(G47), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n558), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AND4_X1   g177(.A1(KEYINPUT78), .A2(new_n596), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n601), .B1(KEYINPUT77), .B2(new_n595), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT78), .B1(new_n604), .B2(new_n598), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n539), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n512), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n525), .A2(G54), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(G171), .ZN(G284));
  OAI21_X1  g192(.A(new_n616), .B1(new_n615), .B2(G171), .ZN(G321));
  AOI21_X1  g193(.A(new_n569), .B1(new_n560), .B2(new_n562), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G286), .B2(G868), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(G297));
  XOR2_X1   g197(.A(new_n621), .B(KEYINPUT80), .Z(G280));
  AND3_X1   g198(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  INV_X1    g201(.A(new_n549), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n615), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n614), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n472), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n465), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n463), .A2(new_n473), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n638), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT13), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT82), .Z(G156));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2438), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT83), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT16), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n649), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n649), .B2(new_n650), .ZN(new_n657));
  OR3_X1    g232(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n656), .B1(new_n654), .B2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n668), .ZN(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n671), .A2(KEYINPUT17), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n671), .B2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n666), .A2(new_n668), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G2100), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT85), .B(G2096), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR3_X1    g258(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n690), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1991), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n703), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n706), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n706), .B2(new_n710), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(G229));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G28), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n715), .B1(new_n717), .B2(new_n720), .C1(new_n636), .C2(new_n718), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n722), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1966), .ZN(new_n725));
  NAND2_X1  g300(.A1(G171), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G5), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n721), .B(new_n725), .C1(G1961), .C2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT95), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n463), .A2(G127), .ZN(new_n731));
  NAND2_X1  g306(.A1(G115), .A2(G2104), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n465), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n473), .A2(G103), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT25), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n733), .B(new_n735), .C1(G139), .C2(new_n472), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n718), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n718), .B2(G33), .ZN(new_n738));
  INV_X1    g313(.A(G2072), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G32), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT26), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G105), .B2(new_n473), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n483), .A2(G129), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n472), .A2(G141), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  AOI21_X1  g325(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n738), .B2(new_n739), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n722), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n549), .B2(new_n722), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1341), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n624), .A2(new_n722), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G4), .B2(new_n722), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n718), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n718), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT29), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n759), .A2(new_n760), .B1(G2090), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n760), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(G2090), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n718), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n718), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n728), .B2(G1961), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n757), .A2(new_n764), .A3(new_n767), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n718), .A2(G26), .ZN(new_n774));
  INV_X1    g349(.A(new_n472), .ZN(new_n775));
  INV_X1    g350(.A(G140), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n775), .A2(KEYINPUT92), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT93), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(G128), .B2(new_n483), .ZN(new_n783));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n775), .B2(new_n776), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n777), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n774), .B1(new_n785), .B2(G29), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n774), .B(new_n786), .S(KEYINPUT28), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2067), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(KEYINPUT24), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n479), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G2084), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n788), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT23), .B1(new_n619), .B2(new_n722), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n722), .A2(G20), .ZN(new_n798));
  MUX2_X1   g373(.A(KEYINPUT23), .B(new_n797), .S(new_n798), .Z(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n730), .A2(new_n773), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G16), .B2(G23), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n804), .B(new_n806), .C1(G16), .C2(G23), .ZN(new_n809));
  INV_X1    g384(.A(G305), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n722), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G6), .B2(new_n722), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT90), .B(KEYINPUT32), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1981), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n808), .B(new_n809), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G22), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G166), .B2(G16), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT91), .B(G1971), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n812), .A2(new_n814), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n722), .A2(G24), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n606), .B2(new_n722), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT89), .B(G1986), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G119), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n482), .A2(KEYINPUT87), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT87), .B1(new_n482), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n472), .A2(G131), .ZN(new_n831));
  OR3_X1    g406(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n465), .A2(G107), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(G2104), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  MUX2_X1   g411(.A(G25), .B(new_n836), .S(G29), .Z(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT35), .B(G1991), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n823), .A2(new_n827), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n802), .B1(new_n842), .B2(new_n843), .ZN(G311));
  INV_X1    g419(.A(G311), .ZN(G150));
  NAND2_X1  g420(.A1(new_n525), .A2(G55), .ZN(new_n846));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n509), .B2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(G651), .A2(new_n849), .B1(new_n539), .B2(G93), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(KEYINPUT96), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT96), .B1(new_n846), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT99), .B(G860), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n846), .A2(new_n850), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n549), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n549), .A2(new_n858), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT97), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n627), .B1(new_n852), .B2(new_n853), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(new_n862), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT98), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT97), .B1(new_n861), .B2(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n865), .A3(new_n862), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n868), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n614), .A2(new_n625), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT38), .B1(new_n868), .B2(new_n872), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n855), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n875), .B1(new_n873), .B2(new_n876), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n857), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT100), .ZN(G145));
  INV_X1    g457(.A(new_n640), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n483), .A2(G130), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n472), .A2(G142), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n465), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n836), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n883), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n640), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT102), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n501), .A2(new_n503), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n497), .A2(new_n498), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n736), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n785), .B(new_n747), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n905), .B(new_n906), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n489), .B(new_n636), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n479), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g494(.A(G166), .B(new_n810), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT78), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n604), .A2(KEYINPUT78), .A3(new_n598), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n924), .A2(G288), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G288), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n803), .B1(new_n603), .B2(new_n605), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(G288), .A3(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n932), .B2(new_n921), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n930), .A2(KEYINPUT104), .A3(new_n931), .A4(new_n920), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n624), .A2(G299), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n614), .A2(new_n619), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT103), .B1(new_n624), .B2(G299), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT41), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n948), .A3(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(new_n629), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n870), .A2(new_n871), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n870), .B2(new_n871), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n947), .B(new_n949), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n953), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n945), .A2(new_n946), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n951), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n940), .B1(new_n935), .B2(new_n939), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n941), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n935), .A2(new_n939), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n854), .A2(new_n615), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n966), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n958), .B1(new_n941), .B2(new_n959), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n961), .A3(new_n964), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n615), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n967), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(KEYINPUT106), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n970), .A2(new_n975), .ZN(G331));
  NAND2_X1  g551(.A1(new_n943), .A2(new_n944), .ZN(new_n977));
  NOR2_X1   g552(.A1(G171), .A2(new_n533), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n575), .B2(G301), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n870), .A3(new_n871), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n870), .B2(new_n871), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT41), .B(new_n977), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(G286), .B2(G171), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n864), .B2(new_n867), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n948), .B1(new_n986), .B2(new_n981), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n956), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n935), .A2(new_n939), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n962), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n947), .B(new_n949), .C1(new_n982), .C2(new_n983), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n956), .A2(new_n981), .A3(new_n986), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n917), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n992), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n996), .ZN(new_n1000));
  AOI21_X1  g575(.A(G37), .B1(new_n1000), .B2(new_n962), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n935), .A2(new_n939), .A3(new_n990), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n990), .B1(new_n935), .B2(new_n939), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT44), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n992), .A2(new_n997), .A3(KEYINPUT43), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n998), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n904), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n466), .A2(new_n474), .A3(new_n478), .A4(G40), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n836), .A2(new_n838), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n836), .A2(new_n838), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2067), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n785), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G1996), .B2(new_n747), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1017), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(G1996), .A3(new_n747), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1986), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n606), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT108), .Z(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1030), .B2(new_n606), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1021), .B(new_n1029), .C1(new_n1033), .C2(new_n1017), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(new_n1039), .C1(new_n1038), .C2(G288), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR3_X1    g617(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT115), .B(G86), .Z(new_n1046));
  OAI21_X1  g621(.A(new_n586), .B1(new_n540), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1037), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT49), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1042), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1037), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(new_n1038), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1041), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n904), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1016), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1015), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1971), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n904), .B2(new_n1012), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1065), .B2(new_n1016), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1067), .A3(KEYINPUT116), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT50), .B(G1384), .C1(new_n902), .C2(new_n903), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT111), .B(G2090), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1062), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G303), .A2(G8), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT55), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1067), .B1(new_n1069), .B2(KEYINPUT110), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1072), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1013), .A2(new_n1081), .A3(KEYINPUT50), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1079), .A2(new_n1059), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1062), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT112), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1062), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1078), .A2(new_n1085), .A3(G8), .A4(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1057), .A2(new_n1077), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1036), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT117), .B(G2084), .Z(new_n1091));
  NAND4_X1  g666(.A1(new_n1079), .A2(new_n1059), .A3(new_n1082), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1060), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1095), .B2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1090), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n1097), .B2(KEYINPUT122), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1036), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(new_n1090), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AND4_X1   g679(.A1(KEYINPUT123), .A2(new_n1100), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1102), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT62), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(KEYINPUT123), .A3(new_n1102), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT124), .B(G1961), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1079), .A2(new_n1059), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1082), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1060), .B2(G2078), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1015), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(KEYINPUT53), .A3(new_n770), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G171), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1108), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT119), .B1(G299), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n619), .A2(new_n1129), .A3(KEYINPUT57), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n619), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT120), .B1(new_n619), .B2(KEYINPUT57), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1128), .A2(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1071), .A2(new_n800), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1121), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n760), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1035), .A2(new_n1022), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n614), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1133), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n624), .A2(KEYINPUT60), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1139), .A2(new_n1140), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1015), .A2(new_n1059), .A3(new_n707), .A4(new_n1058), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1035), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  AOI22_X1  g734(.A1(new_n1157), .A2(KEYINPUT121), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1121), .A2(new_n1161), .A3(new_n707), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1156), .B1(new_n1163), .B2(new_n549), .ZN(new_n1164));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n627), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1152), .B(new_n1155), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1142), .B1(new_n1150), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n474), .A2(KEYINPUT53), .A3(G40), .A4(new_n770), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(G2105), .B2(new_n477), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n1015), .A3(new_n1058), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1118), .A2(new_n1120), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(G301), .B1(new_n1172), .B2(KEYINPUT125), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(KEYINPUT125), .B2(new_n1172), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT54), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1123), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(G301), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1124), .B1(G171), .B2(new_n1172), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1174), .A2(new_n1177), .B1(new_n1178), .B2(new_n1175), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1167), .A2(new_n1168), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1089), .B1(new_n1126), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1085), .A2(G8), .A3(new_n1087), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1076), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1183), .A2(KEYINPUT63), .A3(new_n575), .A4(new_n1101), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1057), .A2(new_n1088), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT118), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1101), .A2(new_n575), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1187), .B1(new_n1089), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1187), .B(new_n1188), .C1(new_n1182), .C2(new_n1076), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT118), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1190), .A2(new_n1191), .A3(new_n1088), .A4(new_n1057), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1186), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1038), .B(new_n803), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1053), .B1(new_n1194), .B2(new_n1045), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1088), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1057), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1034), .B1(new_n1181), .B2(new_n1198), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1032), .A2(new_n1018), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT48), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1029), .A2(new_n1021), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  XOR2_X1   g780(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1017), .B2(new_n707), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n707), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1023), .A2(new_n748), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1207), .B1(new_n1209), .B2(new_n1017), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT47), .ZN(new_n1211));
  OAI22_X1  g786(.A1(new_n1029), .A2(new_n1020), .B1(G2067), .B2(new_n785), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1211), .B1(new_n1017), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1205), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1199), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g790(.A1(new_n684), .A2(G319), .A3(new_n685), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1217), .B1(new_n662), .B2(new_n663), .ZN(new_n1218));
  NOR3_X1   g792(.A1(new_n712), .A2(new_n713), .A3(new_n1218), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n1219), .B(new_n918), .C1(new_n1008), .C2(new_n1009), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


