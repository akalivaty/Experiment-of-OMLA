

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767;

  NAND2_X1 U366 ( .A1(n419), .A2(n433), .ZN(n362) );
  INV_X1 U367 ( .A(n546), .ZN(n367) );
  NAND2_X1 U368 ( .A1(n592), .A2(n590), .ZN(n687) );
  INV_X4 U369 ( .A(G953), .ZN(n759) );
  BUF_X1 U370 ( .A(G104), .Z(n399) );
  NOR2_X2 U371 ( .A1(n585), .A2(n661), .ZN(n587) );
  XNOR2_X2 U372 ( .A(n587), .B(n586), .ZN(n763) );
  NOR2_X2 U373 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U374 ( .A1(n546), .A2(n434), .ZN(n419) );
  XNOR2_X2 U375 ( .A(n549), .B(KEYINPUT1), .ZN(n546) );
  NAND2_X2 U376 ( .A1(n344), .A2(n626), .ZN(n722) );
  NAND2_X2 U377 ( .A1(n407), .A2(n410), .ZN(n344) );
  NAND2_X1 U378 ( .A1(n345), .A2(n361), .ZN(n369) );
  NAND2_X1 U379 ( .A1(n351), .A2(n365), .ZN(n345) );
  AND2_X4 U380 ( .A1(n722), .A2(n723), .ZN(n731) );
  XOR2_X2 U381 ( .A(KEYINPUT15), .B(G902), .Z(n492) );
  NOR2_X2 U382 ( .A1(n633), .A2(n736), .ZN(n636) );
  NOR2_X2 U383 ( .A1(n721), .A2(n736), .ZN(n400) );
  XOR2_X1 U384 ( .A(G119), .B(KEYINPUT68), .Z(n453) );
  BUF_X1 U385 ( .A(G128), .Z(n657) );
  AND2_X1 U386 ( .A1(n380), .A2(KEYINPUT2), .ZN(n346) );
  XOR2_X1 U387 ( .A(KEYINPUT107), .B(KEYINPUT63), .Z(n347) );
  XOR2_X1 U388 ( .A(n643), .B(n642), .Z(n348) );
  XOR2_X1 U389 ( .A(n450), .B(n533), .Z(n349) );
  NAND2_X2 U390 ( .A1(n372), .A2(n349), .ZN(n436) );
  NAND2_X2 U391 ( .A1(n358), .A2(n675), .ZN(n445) );
  AND2_X2 U392 ( .A1(n425), .A2(n448), .ZN(n424) );
  AND2_X2 U393 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X2 U394 ( .A(n368), .B(n540), .ZN(n717) );
  NOR2_X1 U395 ( .A1(n684), .A2(n564), .ZN(n565) );
  XOR2_X2 U396 ( .A(n593), .B(KEYINPUT6), .Z(n601) );
  XNOR2_X2 U397 ( .A(n461), .B(n442), .ZN(n593) );
  NOR2_X1 U398 ( .A1(n679), .A2(n678), .ZN(n588) );
  INV_X1 U399 ( .A(n687), .ZN(n374) );
  NAND2_X1 U400 ( .A1(n687), .A2(n434), .ZN(n433) );
  OR2_X1 U401 ( .A1(n734), .A2(G902), .ZN(n426) );
  AND2_X1 U402 ( .A1(n411), .A2(n756), .ZN(n410) );
  NOR2_X1 U403 ( .A1(n680), .A2(n660), .ZN(n608) );
  NAND2_X1 U404 ( .A1(n375), .A2(n374), .ZN(n579) );
  INV_X1 U405 ( .A(n596), .ZN(n375) );
  NOR2_X1 U406 ( .A1(n687), .A2(n434), .ZN(n388) );
  XNOR2_X2 U407 ( .A(n743), .B(n483), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n428), .B(n427), .ZN(n510) );
  NOR2_X1 U409 ( .A1(n728), .A2(n736), .ZN(n730) );
  INV_X1 U410 ( .A(n740), .ZN(n381) );
  BUF_X1 U411 ( .A(n393), .Z(n740) );
  INV_X1 U412 ( .A(n627), .ZN(n380) );
  XNOR2_X1 U413 ( .A(n377), .B(n376), .ZN(n383) );
  INV_X1 U414 ( .A(n362), .ZN(n418) );
  NOR2_X1 U415 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U416 ( .A1(n367), .A2(n388), .ZN(n417) );
  XNOR2_X1 U417 ( .A(n354), .B(n446), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n382), .B(n718), .ZN(n719) );
  AND2_X1 U419 ( .A1(n388), .A2(n366), .ZN(n360) );
  AND2_X1 U420 ( .A1(n433), .A2(n366), .ZN(n359) );
  AND2_X1 U421 ( .A1(n352), .A2(n534), .ZN(n435) );
  BUF_X1 U422 ( .A(n743), .Z(n396) );
  XNOR2_X1 U423 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U424 ( .A(n744), .B(n534), .ZN(n483) );
  NAND2_X1 U425 ( .A1(G214), .A2(n496), .ZN(n675) );
  INV_X1 U426 ( .A(n492), .ZN(n624) );
  INV_X1 U427 ( .A(n391), .ZN(n376) );
  INV_X1 U428 ( .A(n736), .ZN(n350) );
  INV_X1 U429 ( .A(KEYINPUT2), .ZN(n378) );
  XNOR2_X1 U430 ( .A(KEYINPUT67), .B(G469), .ZN(n385) );
  XOR2_X1 U431 ( .A(G125), .B(G146), .Z(n488) );
  XOR2_X1 U432 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n391) );
  XNOR2_X1 U433 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n480) );
  NAND2_X1 U434 ( .A1(n364), .A2(n417), .ZN(n351) );
  NAND2_X1 U435 ( .A1(n436), .A2(n352), .ZN(n443) );
  NAND2_X1 U436 ( .A1(n394), .A2(n449), .ZN(n352) );
  NAND2_X1 U437 ( .A1(n353), .A2(n558), .ZN(n559) );
  NAND2_X1 U438 ( .A1(n353), .A2(n541), .ZN(n554) );
  NOR2_X2 U439 ( .A1(n564), .A2(n530), .ZN(n354) );
  XNOR2_X2 U440 ( .A(n355), .B(KEYINPUT0), .ZN(n564) );
  NAND2_X1 U441 ( .A1(n607), .A2(n498), .ZN(n355) );
  XNOR2_X2 U442 ( .A(n356), .B(n491), .ZN(n628) );
  XNOR2_X2 U443 ( .A(n357), .B(n482), .ZN(n743) );
  XNOR2_X2 U444 ( .A(n523), .B(n506), .ZN(n357) );
  XNOR2_X1 U445 ( .A(n453), .B(KEYINPUT3), .ZN(n744) );
  INV_X1 U446 ( .A(n358), .ZN(n622) );
  XNOR2_X2 U447 ( .A(n495), .B(n387), .ZN(n358) );
  NAND2_X1 U448 ( .A1(n611), .A2(n358), .ZN(n658) );
  NAND2_X1 U449 ( .A1(n419), .A2(n359), .ZN(n364) );
  NAND2_X1 U450 ( .A1(n360), .A2(n367), .ZN(n365) );
  NAND2_X1 U451 ( .A1(n362), .A2(KEYINPUT101), .ZN(n361) );
  INV_X1 U452 ( .A(KEYINPUT101), .ZN(n366) );
  NAND2_X1 U453 ( .A1(n429), .A2(n431), .ZN(n405) );
  XNOR2_X2 U454 ( .A(n430), .B(n444), .ZN(n429) );
  XNOR2_X1 U455 ( .A(n415), .B(KEYINPUT19), .ZN(n607) );
  NAND2_X1 U456 ( .A1(n536), .A2(n537), .ZN(n368) );
  NAND2_X1 U457 ( .A1(n369), .A2(n601), .ZN(n404) );
  NAND2_X1 U458 ( .A1(n420), .A2(KEYINPUT44), .ZN(n430) );
  XNOR2_X2 U459 ( .A(n569), .B(KEYINPUT35), .ZN(n420) );
  XNOR2_X1 U460 ( .A(n370), .B(n347), .ZN(G57) );
  NAND2_X1 U461 ( .A1(n371), .A2(n350), .ZN(n370) );
  XNOR2_X1 U462 ( .A(n644), .B(n348), .ZN(n371) );
  INV_X1 U463 ( .A(n532), .ZN(n372) );
  XNOR2_X2 U464 ( .A(n373), .B(n582), .ZN(n610) );
  NAND2_X1 U465 ( .A1(n581), .A2(n589), .ZN(n373) );
  NAND2_X1 U466 ( .A1(n431), .A2(n429), .ZN(n377) );
  NAND2_X1 U467 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U468 ( .A1(n346), .A2(n381), .ZN(n723) );
  XNOR2_X1 U469 ( .A(n379), .B(n378), .ZN(n711) );
  INV_X1 U470 ( .A(n423), .ZN(n382) );
  XNOR2_X1 U471 ( .A(n399), .B(G110), .ZN(n533) );
  INV_X1 U472 ( .A(G134), .ZN(n451) );
  NOR2_X1 U473 ( .A1(n624), .A2(KEYINPUT78), .ZN(n412) );
  OR2_X1 U474 ( .A1(G902), .A2(G237), .ZN(n496) );
  INV_X1 U475 ( .A(G472), .ZN(n442) );
  NOR2_X1 U476 ( .A1(G953), .A2(G237), .ZN(n514) );
  NAND2_X1 U477 ( .A1(n423), .A2(n384), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U479 ( .A(KEYINPUT102), .B(KEYINPUT30), .ZN(n440) );
  NAND2_X1 U480 ( .A1(n593), .A2(n675), .ZN(n441) );
  XNOR2_X1 U481 ( .A(G113), .B(G137), .ZN(n457) );
  XNOR2_X1 U482 ( .A(n447), .B(KEYINPUT69), .ZN(n446) );
  INV_X1 U483 ( .A(KEYINPUT22), .ZN(n447) );
  INV_X1 U484 ( .A(n592), .ZN(n555) );
  NOR2_X1 U485 ( .A1(G952), .A2(n759), .ZN(n736) );
  INV_X1 U486 ( .A(KEYINPUT81), .ZN(n444) );
  XNOR2_X1 U487 ( .A(n450), .B(n533), .ZN(n449) );
  XOR2_X1 U488 ( .A(KEYINPUT65), .B(G101), .Z(n534) );
  INV_X1 U489 ( .A(KEYINPUT73), .ZN(n434) );
  XOR2_X1 U490 ( .A(G116), .B(KEYINPUT5), .Z(n455) );
  INV_X1 U491 ( .A(KEYINPUT8), .ZN(n427) );
  NAND2_X1 U492 ( .A1(n759), .A2(G234), .ZN(n428) );
  XNOR2_X1 U493 ( .A(G122), .B(KEYINPUT7), .ZN(n501) );
  XOR2_X1 U494 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n502) );
  XOR2_X1 U495 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n518) );
  XNOR2_X1 U496 ( .A(G143), .B(KEYINPUT94), .ZN(n517) );
  XOR2_X1 U497 ( .A(G140), .B(G131), .Z(n516) );
  NAND2_X1 U498 ( .A1(G237), .A2(G234), .ZN(n474) );
  XNOR2_X1 U499 ( .A(n622), .B(n406), .ZN(n676) );
  XNOR2_X1 U500 ( .A(KEYINPUT38), .B(KEYINPUT72), .ZN(n406) );
  AND2_X2 U501 ( .A1(n439), .A2(n437), .ZN(n756) );
  NOR2_X1 U502 ( .A1(n672), .A2(n438), .ZN(n437) );
  INV_X1 U503 ( .A(n674), .ZN(n438) );
  XOR2_X1 U504 ( .A(G119), .B(KEYINPUT23), .Z(n467) );
  XOR2_X1 U505 ( .A(KEYINPUT41), .B(n588), .Z(n708) );
  INV_X1 U506 ( .A(KEYINPUT33), .ZN(n414) );
  INV_X1 U507 ( .A(KEYINPUT86), .ZN(n493) );
  INV_X1 U508 ( .A(KEYINPUT74), .ZN(n582) );
  XNOR2_X1 U509 ( .A(n630), .B(n629), .ZN(n631) );
  INV_X1 U510 ( .A(n554), .ZN(n401) );
  INV_X1 U511 ( .A(KEYINPUT122), .ZN(n402) );
  NOR2_X1 U512 ( .A1(n385), .A2(G902), .ZN(n384) );
  XOR2_X1 U513 ( .A(G137), .B(G140), .Z(n531) );
  XOR2_X1 U514 ( .A(G143), .B(n657), .Z(n386) );
  XOR2_X1 U515 ( .A(n494), .B(n493), .Z(n387) );
  XOR2_X1 U516 ( .A(n465), .B(n464), .Z(n389) );
  AND2_X1 U517 ( .A1(n689), .A2(n555), .ZN(n390) );
  XNOR2_X1 U518 ( .A(KEYINPUT59), .B(KEYINPUT85), .ZN(n392) );
  NAND2_X1 U519 ( .A1(n766), .A2(n652), .ZN(n561) );
  XNOR2_X1 U520 ( .A(n405), .B(n391), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n751), .B(G146), .ZN(n394) );
  XNOR2_X1 U522 ( .A(n751), .B(G146), .ZN(n395) );
  XNOR2_X1 U523 ( .A(n751), .B(G146), .ZN(n532) );
  XNOR2_X1 U524 ( .A(n404), .B(n414), .ZN(n684) );
  XNOR2_X1 U525 ( .A(n469), .B(n468), .ZN(n470) );
  BUF_X1 U526 ( .A(n549), .Z(n596) );
  BUF_X1 U527 ( .A(n607), .Z(n397) );
  NOR2_X2 U528 ( .A1(n628), .A2(n492), .ZN(n495) );
  BUF_X1 U529 ( .A(n628), .Z(n398) );
  XNOR2_X1 U530 ( .A(n472), .B(n753), .ZN(n734) );
  XNOR2_X1 U531 ( .A(n400), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U532 ( .A1(n401), .A2(n390), .ZN(n652) );
  XNOR2_X2 U533 ( .A(n559), .B(KEYINPUT32), .ZN(n766) );
  XNOR2_X1 U534 ( .A(n403), .B(n402), .ZN(G63) );
  NAND2_X1 U535 ( .A1(n640), .A2(n350), .ZN(n403) );
  XNOR2_X1 U536 ( .A(n617), .B(KEYINPUT48), .ZN(n439) );
  NOR2_X1 U537 ( .A1(n763), .A2(n767), .ZN(n600) );
  NOR2_X2 U538 ( .A1(n601), .A2(n542), .ZN(n645) );
  INV_X1 U539 ( .A(n756), .ZN(n627) );
  NAND2_X1 U540 ( .A1(n624), .A2(KEYINPUT78), .ZN(n408) );
  NAND2_X1 U541 ( .A1(n393), .A2(KEYINPUT78), .ZN(n409) );
  NAND2_X1 U542 ( .A1(n383), .A2(n412), .ZN(n411) );
  NAND2_X1 U543 ( .A1(n418), .A2(n417), .ZN(n562) );
  NOR2_X1 U544 ( .A1(n618), .A2(n415), .ZN(n604) );
  XNOR2_X2 U545 ( .A(n445), .B(n497), .ZN(n415) );
  XNOR2_X2 U546 ( .A(n416), .B(G113), .ZN(n523) );
  XNOR2_X2 U547 ( .A(G122), .B(G104), .ZN(n416) );
  INV_X1 U548 ( .A(n420), .ZN(n421) );
  NAND2_X1 U549 ( .A1(n420), .A2(n570), .ZN(n571) );
  XNOR2_X1 U550 ( .A(n421), .B(G122), .ZN(n765) );
  NAND2_X2 U551 ( .A1(n424), .A2(n422), .ZN(n549) );
  INV_X1 U552 ( .A(n717), .ZN(n423) );
  NAND2_X1 U553 ( .A1(n717), .A2(n385), .ZN(n425) );
  XNOR2_X2 U554 ( .A(n426), .B(n389), .ZN(n592) );
  NAND2_X1 U555 ( .A1(n510), .A2(G221), .ZN(n466) );
  AND2_X2 U556 ( .A1(n432), .A2(n573), .ZN(n431) );
  NAND2_X1 U557 ( .A1(n571), .A2(n572), .ZN(n432) );
  NAND2_X1 U558 ( .A1(n435), .A2(n436), .ZN(n537) );
  XNOR2_X1 U559 ( .A(n441), .B(n440), .ZN(n580) );
  NAND2_X1 U560 ( .A1(n443), .A2(n535), .ZN(n536) );
  NAND2_X1 U561 ( .A1(n385), .A2(G902), .ZN(n448) );
  INV_X1 U562 ( .A(n531), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n727), .B(n726), .ZN(n728) );
  INV_X1 U564 ( .A(KEYINPUT46), .ZN(n599) );
  XNOR2_X1 U565 ( .A(n600), .B(n599), .ZN(n616) );
  BUF_X1 U566 ( .A(n684), .Z(n707) );
  INV_X1 U567 ( .A(KEYINPUT24), .ZN(n468) );
  INV_X1 U568 ( .A(KEYINPUT83), .ZN(n497) );
  XNOR2_X1 U569 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U570 ( .A(n725), .B(n392), .ZN(n726) );
  XNOR2_X1 U571 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X2 U572 ( .A(G143), .B(G128), .ZN(n487) );
  XNOR2_X2 U573 ( .A(n487), .B(n451), .ZN(n504) );
  XNOR2_X1 U574 ( .A(KEYINPUT4), .B(G131), .ZN(n452) );
  XNOR2_X2 U575 ( .A(n504), .B(n452), .ZN(n751) );
  XNOR2_X1 U576 ( .A(n395), .B(n483), .ZN(n460) );
  NAND2_X1 U577 ( .A1(n514), .A2(G210), .ZN(n454) );
  XNOR2_X1 U578 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U579 ( .A(n456), .B(KEYINPUT92), .Z(n458) );
  XNOR2_X1 U580 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U581 ( .A(n460), .B(n459), .ZN(n641) );
  NOR2_X1 U582 ( .A1(G902), .A2(n641), .ZN(n461) );
  XOR2_X1 U583 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n465) );
  NAND2_X1 U584 ( .A1(n624), .A2(G234), .ZN(n463) );
  XNOR2_X1 U585 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n462) );
  XNOR2_X1 U586 ( .A(n463), .B(n462), .ZN(n499) );
  NAND2_X1 U587 ( .A1(G217), .A2(n499), .ZN(n464) );
  XNOR2_X1 U588 ( .A(n488), .B(KEYINPUT10), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n531), .B(n521), .ZN(n753) );
  XNOR2_X1 U590 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U591 ( .A(n657), .B(G110), .ZN(n469) );
  XNOR2_X1 U592 ( .A(KEYINPUT100), .B(n555), .ZN(n691) );
  NOR2_X1 U593 ( .A1(G898), .A2(n759), .ZN(n473) );
  XNOR2_X1 U594 ( .A(KEYINPUT88), .B(n473), .ZN(n747) );
  XNOR2_X1 U595 ( .A(n474), .B(KEYINPUT14), .ZN(n476) );
  NAND2_X1 U596 ( .A1(n476), .A2(G902), .ZN(n475) );
  XNOR2_X1 U597 ( .A(n475), .B(KEYINPUT89), .ZN(n574) );
  NAND2_X1 U598 ( .A1(n747), .A2(n574), .ZN(n479) );
  NAND2_X1 U599 ( .A1(G952), .A2(n476), .ZN(n706) );
  NOR2_X1 U600 ( .A1(G953), .A2(n706), .ZN(n477) );
  XOR2_X1 U601 ( .A(KEYINPUT87), .B(n477), .Z(n577) );
  INV_X1 U602 ( .A(n577), .ZN(n478) );
  NAND2_X1 U603 ( .A1(n479), .A2(n478), .ZN(n498) );
  XOR2_X2 U604 ( .A(G116), .B(G107), .Z(n506) );
  XOR2_X1 U605 ( .A(G110), .B(KEYINPUT16), .Z(n481) );
  XNOR2_X1 U606 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n485) );
  NAND2_X1 U608 ( .A1(G224), .A2(n759), .ZN(n484) );
  XNOR2_X1 U609 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U610 ( .A(n486), .B(KEYINPUT4), .Z(n490) );
  XNOR2_X1 U611 ( .A(n386), .B(n488), .ZN(n489) );
  NAND2_X1 U612 ( .A1(G210), .A2(n496), .ZN(n494) );
  NAND2_X1 U613 ( .A1(n499), .A2(G221), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n500), .B(KEYINPUT21), .ZN(n692) );
  XNOR2_X1 U615 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U616 ( .A(n503), .B(KEYINPUT9), .Z(n509) );
  BUF_X1 U617 ( .A(n504), .Z(n505) );
  INV_X1 U618 ( .A(n505), .ZN(n507) );
  XNOR2_X1 U619 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U620 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U621 ( .A1(n510), .A2(G217), .ZN(n511) );
  XNOR2_X1 U622 ( .A(n512), .B(n511), .ZN(n637) );
  NOR2_X1 U623 ( .A1(n637), .A2(G902), .ZN(n513) );
  XOR2_X1 U624 ( .A(G478), .B(n513), .Z(n543) );
  INV_X1 U625 ( .A(n543), .ZN(n567) );
  XNOR2_X1 U626 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n527) );
  NAND2_X1 U627 ( .A1(n514), .A2(G214), .ZN(n515) );
  XNOR2_X1 U628 ( .A(n516), .B(n515), .ZN(n520) );
  XNOR2_X1 U629 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U630 ( .A(n520), .B(n519), .Z(n525) );
  INV_X1 U631 ( .A(n521), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n525), .B(n524), .ZN(n725) );
  NOR2_X1 U634 ( .A1(G902), .A2(n725), .ZN(n526) );
  XNOR2_X1 U635 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U636 ( .A(G475), .B(n528), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n678) );
  NOR2_X1 U638 ( .A1(n692), .A2(n678), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n529), .B(KEYINPUT99), .ZN(n530) );
  INV_X1 U640 ( .A(n534), .ZN(n535) );
  NAND2_X1 U641 ( .A1(G227), .A2(n759), .ZN(n539) );
  XNOR2_X1 U642 ( .A(G107), .B(KEYINPUT75), .ZN(n538) );
  BUF_X1 U643 ( .A(n546), .Z(n541) );
  INV_X1 U644 ( .A(n541), .ZN(n619) );
  OR2_X1 U645 ( .A1(n691), .A2(n554), .ZN(n542) );
  NAND2_X1 U646 ( .A1(n543), .A2(n566), .ZN(n653) );
  INV_X1 U647 ( .A(n653), .ZN(n666) );
  INV_X1 U648 ( .A(n566), .ZN(n544) );
  NAND2_X1 U649 ( .A1(n544), .A2(n567), .ZN(n661) );
  INV_X1 U650 ( .A(n661), .ZN(n663) );
  NOR2_X1 U651 ( .A1(n666), .A2(n663), .ZN(n545) );
  XNOR2_X1 U652 ( .A(n545), .B(KEYINPUT98), .ZN(n680) );
  INV_X1 U653 ( .A(n564), .ZN(n547) );
  INV_X1 U654 ( .A(n593), .ZN(n689) );
  INV_X1 U655 ( .A(n692), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n689), .A2(n562), .ZN(n699) );
  NAND2_X1 U657 ( .A1(n547), .A2(n699), .ZN(n548) );
  XNOR2_X1 U658 ( .A(n548), .B(KEYINPUT31), .ZN(n667) );
  NOR2_X1 U659 ( .A1(n564), .A2(n579), .ZN(n550) );
  NAND2_X1 U660 ( .A1(n550), .A2(n689), .ZN(n551) );
  XNOR2_X1 U661 ( .A(KEYINPUT93), .B(n551), .ZN(n647) );
  NOR2_X1 U662 ( .A1(n667), .A2(n647), .ZN(n552) );
  NOR2_X1 U663 ( .A1(n680), .A2(n552), .ZN(n553) );
  NOR2_X1 U664 ( .A1(n645), .A2(n553), .ZN(n573) );
  INV_X1 U665 ( .A(n601), .ZN(n563) );
  NAND2_X1 U666 ( .A1(n563), .A2(n691), .ZN(n556) );
  NOR2_X1 U667 ( .A1(n541), .A2(n556), .ZN(n557) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n557), .ZN(n558) );
  INV_X1 U669 ( .A(KEYINPUT44), .ZN(n570) );
  NAND2_X1 U670 ( .A1(KEYINPUT82), .A2(n570), .ZN(n560) );
  XNOR2_X1 U671 ( .A(n561), .B(n560), .ZN(n572) );
  XNOR2_X1 U672 ( .A(n565), .B(KEYINPUT34), .ZN(n568) );
  NOR2_X1 U673 ( .A1(n567), .A2(n566), .ZN(n609) );
  NAND2_X1 U674 ( .A1(n568), .A2(n609), .ZN(n569) );
  XOR2_X1 U675 ( .A(KEYINPUT80), .B(KEYINPUT39), .Z(n584) );
  NAND2_X1 U676 ( .A1(G953), .A2(n574), .ZN(n575) );
  NOR2_X1 U677 ( .A1(G900), .A2(n575), .ZN(n576) );
  NOR2_X1 U678 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U679 ( .A(KEYINPUT77), .B(n578), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n610), .A2(n676), .ZN(n583) );
  XNOR2_X1 U681 ( .A(n583), .B(n584), .ZN(n585) );
  NOR2_X1 U682 ( .A1(n585), .A2(n653), .ZN(n672) );
  XNOR2_X1 U683 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n586) );
  NAND2_X1 U684 ( .A1(n676), .A2(n675), .ZN(n679) );
  XOR2_X1 U685 ( .A(KEYINPUT103), .B(KEYINPUT28), .Z(n595) );
  NAND2_X1 U686 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U687 ( .A1(n592), .A2(n591), .ZN(n602) );
  NAND2_X1 U688 ( .A1(n593), .A2(n602), .ZN(n594) );
  XNOR2_X1 U689 ( .A(n595), .B(n594), .ZN(n597) );
  NOR2_X1 U690 ( .A1(n597), .A2(n596), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n708), .A2(n606), .ZN(n598) );
  XOR2_X1 U692 ( .A(KEYINPUT42), .B(n598), .Z(n767) );
  AND2_X1 U693 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U694 ( .A1(n663), .A2(n603), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT36), .B(n604), .Z(n605) );
  NOR2_X1 U696 ( .A1(n541), .A2(n605), .ZN(n669) );
  NAND2_X1 U697 ( .A1(n397), .A2(n606), .ZN(n660) );
  XNOR2_X1 U698 ( .A(n608), .B(KEYINPUT47), .ZN(n612) );
  AND2_X1 U699 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n612), .A2(n658), .ZN(n613) );
  NOR2_X1 U701 ( .A1(n669), .A2(n613), .ZN(n614) );
  XOR2_X1 U702 ( .A(KEYINPUT66), .B(n614), .Z(n615) );
  NOR2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n620), .A2(n675), .ZN(n621) );
  XNOR2_X1 U705 ( .A(KEYINPUT43), .B(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n674) );
  XNOR2_X1 U707 ( .A(n624), .B(KEYINPUT79), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n625), .A2(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n731), .A2(G210), .ZN(n632) );
  XOR2_X1 U710 ( .A(KEYINPUT84), .B(KEYINPUT55), .Z(n630) );
  XNOR2_X1 U711 ( .A(n398), .B(KEYINPUT54), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U713 ( .A(KEYINPUT119), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT56), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n636), .B(n635), .ZN(G51) );
  NAND2_X1 U716 ( .A1(n731), .A2(G478), .ZN(n639) );
  INV_X1 U717 ( .A(n637), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U719 ( .A(KEYINPUT105), .B(KEYINPUT62), .Z(n643) );
  XNOR2_X1 U720 ( .A(n641), .B(KEYINPUT106), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n731), .A2(G472), .ZN(n644) );
  XOR2_X1 U722 ( .A(G101), .B(n645), .Z(G3) );
  NAND2_X1 U723 ( .A1(n647), .A2(n663), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(n399), .ZN(G6) );
  XNOR2_X1 U725 ( .A(G107), .B(KEYINPUT27), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT26), .B(KEYINPUT108), .Z(n649) );
  NAND2_X1 U727 ( .A1(n647), .A2(n666), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(G9) );
  XNOR2_X1 U730 ( .A(G110), .B(n652), .ZN(G12) );
  NOR2_X1 U731 ( .A1(n653), .A2(n660), .ZN(n655) );
  XNOR2_X1 U732 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U734 ( .A(n657), .B(n656), .Z(G30) );
  XNOR2_X1 U735 ( .A(G143), .B(KEYINPUT110), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(G45) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U738 ( .A(G146), .B(n662), .Z(G48) );
  XOR2_X1 U739 ( .A(G113), .B(KEYINPUT111), .Z(n665) );
  NAND2_X1 U740 ( .A1(n667), .A2(n663), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n665), .B(n664), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U743 ( .A(n668), .B(G116), .ZN(G18) );
  XNOR2_X1 U744 ( .A(n669), .B(KEYINPUT112), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(KEYINPUT37), .ZN(n671) );
  XNOR2_X1 U746 ( .A(G125), .B(n671), .ZN(G27) );
  XNOR2_X1 U747 ( .A(G134), .B(n672), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(KEYINPUT113), .ZN(G36) );
  XNOR2_X1 U749 ( .A(G140), .B(n674), .ZN(G42) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n716) );
  NOR2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n683) );
  NOR2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n681), .B(KEYINPUT116), .ZN(n682) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U756 ( .A1(n685), .A2(n707), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n686), .B(KEYINPUT117), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n541), .A2(n687), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT50), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n697) );
  XOR2_X1 U761 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n694) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(KEYINPUT114), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n701), .A2(n708), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U770 ( .A(KEYINPUT52), .B(n704), .Z(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n713) );
  INV_X1 U772 ( .A(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n714), .A2(n759), .ZN(n715) );
  XNOR2_X1 U777 ( .A(n716), .B(n715), .ZN(G75) );
  NAND2_X1 U778 ( .A1(n731), .A2(G469), .ZN(n720) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n718) );
  AND2_X1 U780 ( .A1(G475), .A2(n723), .ZN(n724) );
  NAND2_X1 U781 ( .A1(n722), .A2(n724), .ZN(n727) );
  XOR2_X1 U782 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n729) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(G60) );
  BUF_X1 U784 ( .A(n731), .Z(n732) );
  NAND2_X1 U785 ( .A1(G217), .A2(n732), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(G66) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n738), .A2(G898), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n739), .B(KEYINPUT123), .ZN(n742) );
  NOR2_X1 U792 ( .A1(G953), .A2(n740), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n749) );
  XNOR2_X1 U794 ( .A(n396), .B(G101), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U796 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U797 ( .A(n749), .B(n748), .Z(n750) );
  XNOR2_X1 U798 ( .A(KEYINPUT124), .B(n750), .ZN(G69) );
  BUF_X1 U799 ( .A(n751), .Z(n752) );
  XNOR2_X1 U800 ( .A(n753), .B(n752), .ZN(n757) );
  XNOR2_X1 U801 ( .A(G227), .B(n757), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(G900), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(G953), .ZN(n762) );
  XNOR2_X1 U804 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n758), .B(KEYINPUT125), .ZN(n760) );
  NAND2_X1 U806 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U807 ( .A1(n762), .A2(n761), .ZN(G72) );
  XNOR2_X1 U808 ( .A(n763), .B(G131), .ZN(n764) );
  XNOR2_X1 U809 ( .A(n764), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U810 ( .A(KEYINPUT126), .B(n765), .ZN(G24) );
  XNOR2_X1 U811 ( .A(n766), .B(G119), .ZN(G21) );
  XOR2_X1 U812 ( .A(G137), .B(n767), .Z(G39) );
endmodule

