//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n193), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n206), .A2(new_n200), .A3(new_n202), .A4(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT0), .B(G128), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n220), .A2(new_n210), .A3(new_n212), .A4(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n210), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n215), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n221), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n199), .A2(G137), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n201), .A2(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n207), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n197), .B(new_n219), .C1(new_n237), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G237), .ZN(new_n243));
  INV_X1    g057(.A(G953), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G210), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT27), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G101), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n219), .A2(KEYINPUT30), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n237), .B2(new_n241), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n221), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n231), .A2(KEYINPUT68), .A3(new_n232), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n231), .B2(new_n232), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n241), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT69), .A3(new_n251), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n207), .A2(new_n263), .A3(new_n240), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n207), .B2(new_n240), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n219), .B1(new_n237), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n197), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI211_X1 g083(.A(KEYINPUT31), .B(new_n249), .C1(new_n262), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n268), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n253), .B(new_n250), .C1(new_n258), .C2(new_n259), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT69), .B1(new_n260), .B2(new_n251), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n196), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n249), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n248), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n219), .B1(new_n237), .B2(new_n241), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n196), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n217), .B1(new_n205), .B2(new_n207), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n258), .B2(new_n259), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n267), .A2(new_n196), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n242), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n279), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n264), .A2(new_n265), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n283), .B1(new_n258), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n196), .B1(new_n293), .B2(KEYINPUT30), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n254), .B2(new_n261), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT31), .B1(new_n295), .B2(new_n249), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n275), .A2(new_n271), .A3(new_n276), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n290), .A3(KEYINPUT71), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n280), .A2(new_n196), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n304), .B2(new_n242), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n286), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n248), .A2(KEYINPUT29), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n275), .A2(new_n242), .A3(new_n279), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n248), .B1(new_n286), .B2(new_n289), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G472), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n187), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n290), .A3(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n316), .B2(new_n298), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT32), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n302), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G210), .B1(G237), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G104), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n322), .B2(G107), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT78), .B1(new_n322), .B2(G107), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(G107), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G104), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n330));
  OR2_X1    g144(.A1(KEYINPUT77), .A2(G107), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT77), .A2(G107), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT78), .A4(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n328), .A2(new_n329), .A3(G101), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT77), .A2(G107), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT77), .A2(G107), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n327), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n323), .A2(new_n324), .ZN(new_n340));
  OAI211_X1 g154(.A(G101), .B(new_n333), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n334), .A2(new_n335), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n196), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G101), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n322), .B1(new_n337), .B2(new_n338), .ZN(new_n349));
  INV_X1    g163(.A(G107), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G104), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n342), .B2(new_n343), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G113), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n194), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n347), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n357), .A2(new_n364), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n194), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n353), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n362), .B(KEYINPUT8), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n369), .B(new_n370), .C1(new_n353), .C2(new_n359), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT73), .B(G125), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n258), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT73), .B(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n218), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n244), .A2(G224), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n373), .A2(new_n375), .B1(KEYINPUT7), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n378), .B(new_n379), .C1(new_n258), .C2(new_n372), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n363), .B(new_n371), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT89), .A3(new_n303), .ZN(new_n382));
  INV_X1    g196(.A(new_n362), .ZN(new_n383));
  INV_X1    g197(.A(new_n343), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n328), .B2(new_n333), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n341), .A2(new_n385), .B1(new_n334), .B2(new_n335), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n334), .A2(new_n335), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n197), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n383), .B1(new_n388), .B2(new_n360), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n363), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n375), .B1(new_n237), .B2(new_n374), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n376), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n383), .C1(new_n388), .C2(new_n360), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n382), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT89), .B1(new_n381), .B2(new_n303), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n321), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n381), .A2(new_n303), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT89), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(new_n320), .A3(new_n395), .A4(new_n382), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G214), .B1(G237), .B2(G902), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT87), .Z(new_n405));
  AND2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G475), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n243), .A2(new_n244), .A3(G214), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(KEYINPUT90), .B2(new_n211), .ZN(new_n410));
  NOR2_X1   g224(.A1(KEYINPUT91), .A2(G143), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT91), .B1(new_n413), .B2(G143), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n243), .A2(new_n244), .A3(G214), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n418));
  INV_X1    g232(.A(G131), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n412), .A2(KEYINPUT18), .A3(G131), .A4(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(G125), .A2(G140), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n374), .B2(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G146), .ZN(new_n425));
  XNOR2_X1  g239(.A(G125), .B(G140), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n209), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT16), .ZN(new_n430));
  INV_X1    g244(.A(G140), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n374), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n424), .B2(new_n430), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n209), .ZN(new_n434));
  OAI211_X1 g248(.A(G146), .B(new_n432), .C1(new_n424), .C2(new_n430), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n206), .B1(new_n412), .B2(new_n416), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n434), .A2(new_n437), .A3(KEYINPUT93), .A4(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n412), .A2(new_n206), .A3(new_n416), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OR3_X1    g257(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n429), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n322), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n438), .A2(new_n439), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n444), .A3(new_n441), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n448), .A3(new_n429), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n448), .B1(new_n453), .B2(new_n429), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n456), .B2(KEYINPUT95), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n407), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n435), .B1(new_n443), .B2(new_n436), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n424), .A2(KEYINPUT19), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n426), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT92), .B1(new_n464), .B2(G146), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n461), .A2(new_n466), .A3(new_n209), .A4(new_n463), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n460), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n429), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n449), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT20), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n454), .B2(new_n470), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n473), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT98), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n190), .A2(G122), .ZN(new_n482));
  INV_X1    g296(.A(G122), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G116), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(new_n325), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n325), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n482), .A2(new_n484), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n331), .A3(new_n332), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n325), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT96), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n227), .A2(new_n229), .A3(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n211), .A2(G128), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n199), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(new_n199), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n488), .A2(new_n492), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n485), .A2(KEYINPUT14), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT14), .ZN(new_n502));
  OAI21_X1  g316(.A(G107), .B1(new_n482), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n493), .A2(new_n199), .A3(new_n494), .ZN(new_n504));
  OAI221_X1 g318(.A(new_n490), .B1(new_n501), .B2(new_n503), .C1(new_n504), .C2(new_n495), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT9), .B(G234), .ZN(new_n506));
  INV_X1    g320(.A(G217), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n506), .A2(new_n507), .A3(G953), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n500), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n500), .B2(new_n505), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n480), .B(new_n303), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT97), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n479), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  OAI211_X1 g328(.A(KEYINPUT97), .B(new_n303), .C1(new_n509), .C2(new_n510), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n516), .B2(new_n479), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT99), .B(G952), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G953), .ZN(new_n519));
  NAND2_X1  g333(.A1(G234), .A2(G237), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n520), .A2(G902), .A3(G953), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT100), .Z(new_n526));
  AND4_X1   g340(.A1(new_n459), .A2(new_n477), .A3(new_n517), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n507), .B1(G234), .B2(new_n303), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n435), .A2(new_n427), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT72), .B(KEYINPUT23), .Z(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n188), .B2(G128), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n188), .A2(G128), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT23), .A4(G119), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G110), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n230), .B2(new_n188), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT74), .B1(new_n534), .B2(new_n535), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n434), .A2(new_n435), .ZN(new_n543));
  OAI221_X1 g357(.A(new_n543), .B1(new_n535), .B2(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n244), .A2(G221), .A3(G234), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT75), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT22), .B(G137), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n545), .B(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n550), .A2(KEYINPUT25), .A3(new_n303), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT25), .B1(new_n550), .B2(new_n303), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n528), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n528), .A2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n319), .A2(new_n406), .A3(new_n527), .A4(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G469), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n222), .A2(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n221), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n353), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT82), .B(new_n563), .C1(new_n258), .C2(new_n353), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n237), .A2(new_n565), .A3(new_n354), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(KEYINPUT12), .A3(new_n566), .A4(new_n208), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT83), .ZN(new_n568));
  INV_X1    g382(.A(new_n208), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n258), .A2(new_n353), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n565), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT83), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT12), .A4(new_n564), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n574));
  INV_X1    g388(.A(new_n564), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n208), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n568), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n385), .A2(new_n579), .A3(new_n352), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n580), .A2(new_n258), .B1(new_n563), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n218), .B1(new_n345), .B2(new_n346), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n569), .ZN(new_n585));
  XNOR2_X1  g399(.A(G110), .B(G140), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n244), .A2(G227), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n578), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n258), .A2(new_n580), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n563), .A2(new_n582), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n217), .B1(new_n386), .B2(new_n387), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n208), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT84), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n583), .A2(new_n584), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(KEYINPUT84), .A3(new_n208), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n601), .B2(new_n585), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n559), .B(new_n303), .C1(new_n591), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT85), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT84), .B1(new_n599), .B2(new_n208), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n597), .B(new_n569), .C1(new_n583), .C2(new_n584), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n585), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n588), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n578), .A2(new_n590), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT85), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n559), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n589), .B1(new_n578), .B2(new_n585), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n601), .A2(new_n590), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n303), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n604), .A2(new_n612), .B1(G469), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G221), .B1(new_n506), .B2(G902), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT76), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT86), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(G469), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n611), .B1(new_n610), .B2(new_n559), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n607), .A2(new_n588), .B1(new_n578), .B2(new_n590), .ZN(new_n622));
  NOR4_X1   g436(.A1(new_n622), .A2(KEYINPUT85), .A3(G469), .A4(G902), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT86), .ZN(new_n625));
  INV_X1    g439(.A(new_n618), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n558), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n343), .B(KEYINPUT101), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT102), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G3));
  OAI21_X1  g446(.A(new_n303), .B1(new_n291), .B2(new_n299), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n317), .B1(new_n633), .B2(G472), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n619), .A2(new_n627), .A3(new_n557), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n477), .A2(new_n459), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n478), .B(new_n303), .C1(new_n509), .C2(new_n510), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n478), .A2(new_n303), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n509), .A2(new_n510), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT33), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n638), .B(new_n639), .C1(new_n641), .C2(G478), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n404), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n398), .B2(new_n402), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n526), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n635), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n471), .B2(new_n474), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT20), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n475), .B(new_n654), .C1(new_n454), .C2(new_n470), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n656), .A2(new_n458), .A3(new_n517), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n645), .A2(new_n650), .A3(new_n526), .A4(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n403), .A2(new_n657), .A3(new_n404), .A4(new_n526), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT104), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n635), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  INV_X1    g477(.A(new_n549), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n545), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n554), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n553), .A2(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n527), .A2(new_n406), .A3(new_n668), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n619), .A2(new_n669), .A3(new_n627), .A4(new_n634), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND3_X1  g486(.A1(new_n520), .A2(G902), .A3(G953), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n521), .B1(G900), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n657), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n675), .A2(new_n645), .A3(new_n668), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n319), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n619), .A4(new_n627), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n619), .A2(new_n627), .A3(new_n319), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT105), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(new_n628), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n674), .B(KEYINPUT39), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n317), .B(new_n301), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n275), .A2(new_n242), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n248), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n304), .A2(new_n242), .A3(new_n279), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n303), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n668), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n403), .B(KEYINPUT38), .Z(new_n697));
  INV_X1    g511(.A(new_n517), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n636), .A2(new_n404), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n687), .A2(new_n688), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  AND3_X1   g517(.A1(new_n636), .A2(new_n642), .A3(new_n674), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n319), .A2(new_n645), .A3(new_n668), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n684), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n622), .B2(G902), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n626), .B(new_n709), .C1(new_n621), .C2(new_n623), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n610), .A2(new_n559), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n604), .B2(new_n612), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT107), .B1(new_n714), .B2(new_n626), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n708), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n646), .A2(new_n643), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n319), .A2(new_n557), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n710), .A2(new_n711), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n714), .A2(KEYINPUT107), .A3(new_n626), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n716), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND2_X1  g538(.A1(new_n660), .A2(new_n658), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(new_n319), .A3(new_n557), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n716), .A2(new_n726), .A3(new_n721), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n712), .A2(new_n715), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n668), .A2(new_n645), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n527), .A3(new_n319), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  INV_X1    g546(.A(new_n403), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n699), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n526), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n633), .A2(G472), .ZN(new_n736));
  INV_X1    g550(.A(new_n278), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n306), .A2(new_n279), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n187), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n557), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n716), .A2(new_n741), .A3(new_n721), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n716), .A2(new_n741), .A3(new_n744), .A4(new_n721), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND3_X1  g561(.A1(new_n719), .A2(new_n720), .A3(new_n645), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n704), .A2(new_n736), .A3(new_n668), .A4(new_n739), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(G125), .Z(G27));
  NOR2_X1   g565(.A1(new_n403), .A2(new_n644), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n624), .A2(new_n626), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n704), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n312), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n300), .A2(KEYINPUT111), .A3(new_n301), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n317), .B2(KEYINPUT32), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n318), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n758), .A2(new_n760), .A3(new_n762), .A4(new_n318), .ZN(new_n765));
  AOI211_X1 g579(.A(KEYINPUT112), .B(new_n556), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT111), .B1(new_n300), .B2(new_n301), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n317), .A2(new_n759), .A3(KEYINPUT32), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n312), .A3(new_n765), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n767), .B1(new_n771), .B2(new_n557), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n756), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n319), .A2(new_n557), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n753), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n704), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n755), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  NAND4_X1  g594(.A1(new_n776), .A2(new_n319), .A3(new_n557), .A4(new_n675), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  INV_X1    g596(.A(new_n752), .ZN(new_n783));
  INV_X1    g597(.A(new_n636), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n642), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT43), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n634), .B1(new_n553), .B2(new_n667), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n613), .A2(new_n614), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT45), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n793), .B2(KEYINPUT45), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(G469), .A2(G902), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT46), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n612), .B2(new_n604), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n797), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n618), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n685), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n792), .B(new_n802), .C1(new_n791), .C2(new_n790), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  XNOR2_X1  g618(.A(new_n801), .B(KEYINPUT47), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n319), .A2(new_n754), .A3(new_n557), .A4(new_n783), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  INV_X1    g622(.A(new_n785), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n626), .A3(new_n405), .A4(new_n557), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT114), .Z(new_n811));
  NAND2_X1  g625(.A1(new_n689), .A2(new_n695), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n714), .B(KEYINPUT49), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n813), .A3(new_n697), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n727), .A2(new_n722), .A3(new_n731), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n743), .B2(new_n745), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n643), .B1(new_n636), .B2(new_n517), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n406), .A3(new_n526), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n635), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n558), .A2(new_n628), .ZN(new_n823));
  INV_X1    g637(.A(new_n670), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n736), .A2(new_n668), .A3(new_n739), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n776), .A2(new_n826), .A3(new_n828), .A4(new_n704), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT116), .B1(new_n749), .B2(new_n753), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n752), .A2(new_n668), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n517), .A2(new_n674), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n656), .A3(new_n458), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n619), .A3(new_n627), .A4(new_n319), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n781), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n825), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n819), .A2(new_n779), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n750), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n626), .A2(new_n734), .A3(new_n624), .A4(new_n674), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n684), .A2(new_n705), .B1(new_n843), .B2(new_n696), .ZN(new_n844));
  AND4_X1   g658(.A1(KEYINPUT52), .A2(new_n682), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n750), .B1(new_n679), .B2(new_n681), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(new_n846), .B2(new_n844), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n817), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n629), .A2(new_n670), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n781), .A2(new_n838), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n822), .A4(new_n831), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n778), .B2(new_n773), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n682), .A2(new_n844), .A3(new_n842), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n844), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT53), .A4(new_n819), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n816), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n858), .A3(new_n819), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT117), .B1(new_n861), .B2(new_n817), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT54), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n849), .A2(new_n859), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n786), .A2(new_n521), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n740), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n644), .A3(new_n697), .A4(new_n729), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT50), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n729), .A2(new_n752), .ZN(new_n876));
  OR4_X1    g690(.A1(new_n521), .A2(new_n876), .A3(new_n556), .A4(new_n812), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n636), .A3(new_n642), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n872), .A2(new_n876), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n828), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n752), .ZN(new_n882));
  INV_X1    g696(.A(new_n805), .ZN(new_n883));
  INV_X1    g697(.A(new_n714), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n626), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT51), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n875), .B(KEYINPUT120), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n880), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n885), .B1(new_n883), .B2(KEYINPUT119), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n882), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n888), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n766), .A2(new_n772), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n879), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT48), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n873), .A2(new_n645), .A3(new_n729), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n519), .C1(new_n877), .C2(new_n643), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n870), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(G952), .A2(G953), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n815), .B1(new_n902), .B2(new_n903), .ZN(G75));
  AOI21_X1  g718(.A(new_n303), .B1(new_n849), .B2(new_n859), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n390), .A2(new_n394), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n392), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n244), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n864), .B(KEYINPUT54), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n797), .B(KEYINPUT57), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n602), .B2(new_n591), .ZN(new_n917));
  INV_X1    g731(.A(new_n796), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n912), .B1(new_n917), .B2(new_n919), .ZN(G54));
  AND3_X1   g734(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(new_n471), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n471), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n912), .ZN(G60));
  AND3_X1   g738(.A1(new_n863), .A2(new_n868), .A3(new_n865), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n868), .B1(new_n863), .B2(new_n865), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n639), .B(KEYINPUT59), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n641), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT121), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n641), .C1(new_n870), .C2(new_n927), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n641), .A2(new_n927), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n912), .B1(new_n914), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n930), .A2(new_n932), .A3(new_n937), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n849), .B2(new_n859), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n912), .B1(new_n942), .B2(new_n666), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n550), .B(KEYINPUT123), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT61), .Z(G66));
  INV_X1    g760(.A(new_n523), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n244), .B1(new_n947), .B2(G224), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n819), .A2(new_n822), .A3(new_n850), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n244), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n907), .B1(G898), .B2(new_n244), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(G69));
  NAND2_X1  g766(.A1(new_n262), .A2(new_n272), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n464), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n803), .A2(new_n807), .A3(new_n781), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n896), .A2(new_n802), .A3(new_n734), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n846), .A2(new_n706), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n955), .A2(new_n779), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n244), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n244), .A2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n954), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n702), .A2(new_n958), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n820), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n783), .B1(new_n820), .B2(new_n966), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n775), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n803), .B(new_n807), .C1(new_n686), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT124), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n965), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n963), .B1(new_n975), .B2(new_n954), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n244), .B1(G227), .B2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n959), .B2(new_n949), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n690), .A2(new_n248), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n912), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n980), .ZN(new_n984));
  INV_X1    g798(.A(new_n949), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n983), .B1(new_n986), .B2(new_n691), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n692), .A2(new_n982), .A3(new_n984), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n860), .B2(new_n862), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT127), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(new_n990), .ZN(G57));
endmodule


