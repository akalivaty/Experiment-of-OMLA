

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U557 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U558 ( .A1(n621), .A2(n734), .ZN(n637) );
  BUF_X1 U559 ( .A(n637), .Z(n677) );
  INV_X1 U560 ( .A(n931), .ZN(n696) );
  NAND2_X1 U561 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U562 ( .A1(G8), .A2(n677), .ZN(n709) );
  NOR2_X1 U563 ( .A1(n642), .A2(n927), .ZN(n635) );
  NOR2_X1 U564 ( .A1(n709), .A2(n696), .ZN(n697) );
  XNOR2_X1 U565 ( .A(n527), .B(KEYINPUT64), .ZN(n547) );
  AND2_X1 U566 ( .A1(G2104), .A2(n529), .ZN(n527) );
  OR2_X1 U567 ( .A1(n709), .A2(n700), .ZN(n523) );
  AND2_X1 U568 ( .A1(n698), .A2(n697), .ZN(n524) );
  XOR2_X1 U569 ( .A(n669), .B(n668), .Z(n525) );
  AND2_X1 U570 ( .A1(n981), .A2(n765), .ZN(n526) );
  NOR2_X1 U571 ( .A1(n689), .A2(n686), .ZN(n667) );
  INV_X1 U572 ( .A(KEYINPUT29), .ZN(n656) );
  AND2_X1 U573 ( .A1(G160), .A2(G40), .ZN(n621) );
  XNOR2_X1 U574 ( .A(n694), .B(KEYINPUT106), .ZN(n705) );
  INV_X1 U575 ( .A(KEYINPUT66), .ZN(n534) );
  NAND2_X1 U576 ( .A1(n523), .A2(n943), .ZN(n701) );
  XNOR2_X1 U577 ( .A(n534), .B(KEYINPUT17), .ZN(n535) );
  XNOR2_X1 U578 ( .A(n536), .B(n535), .ZN(n542) );
  OR2_X1 U579 ( .A1(n753), .A2(n526), .ZN(n754) );
  INV_X1 U580 ( .A(KEYINPUT83), .ZN(n543) );
  NOR2_X1 U581 ( .A1(G651), .A2(n591), .ZN(n796) );
  XNOR2_X1 U582 ( .A(n544), .B(n543), .ZN(n546) );
  INV_X1 U583 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U584 ( .A1(G101), .A2(n547), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n528), .Z(n531) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n529), .ZN(n885) );
  NAND2_X1 U587 ( .A1(n885), .A2(G125), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U589 ( .A(KEYINPUT65), .ZN(n532) );
  XNOR2_X1 U590 ( .A(n533), .B(n532), .ZN(n541) );
  AND2_X1 U591 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U592 ( .A1(G113), .A2(n886), .ZN(n539) );
  NOR2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  INV_X1 U594 ( .A(n542), .ZN(n537) );
  INV_X1 U595 ( .A(n537), .ZN(n882) );
  NAND2_X1 U596 ( .A1(G137), .A2(n882), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X2 U598 ( .A1(n541), .A2(n540), .ZN(G160) );
  NAND2_X1 U599 ( .A1(G138), .A2(n542), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n886), .A2(G114), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n885), .A2(G126), .ZN(n550) );
  INV_X1 U603 ( .A(n547), .ZN(n548) );
  INV_X1 U604 ( .A(n548), .ZN(n881) );
  NAND2_X1 U605 ( .A1(G102), .A2(n881), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G164) );
  XNOR2_X1 U608 ( .A(G543), .B(KEYINPUT0), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT67), .ZN(n591) );
  NAND2_X1 U610 ( .A1(G53), .A2(n796), .ZN(n556) );
  XOR2_X1 U611 ( .A(KEYINPUT68), .B(G651), .Z(n557) );
  NOR2_X1 U612 ( .A1(G543), .A2(n557), .ZN(n554) );
  XOR2_X2 U613 ( .A(KEYINPUT1), .B(n554), .Z(n797) );
  NAND2_X1 U614 ( .A1(G65), .A2(n797), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n561) );
  NOR2_X1 U616 ( .A1(G543), .A2(G651), .ZN(n792) );
  NAND2_X1 U617 ( .A1(n792), .A2(G91), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n591), .A2(n557), .ZN(n793) );
  NAND2_X1 U619 ( .A1(G78), .A2(n793), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U623 ( .A1(G52), .A2(n796), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G64), .A2(n797), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n792), .A2(G90), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G77), .A2(n793), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U630 ( .A1(n569), .A2(n568), .ZN(G171) );
  XNOR2_X1 U631 ( .A(KEYINPUT72), .B(KEYINPUT6), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G51), .A2(n796), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G63), .A2(n797), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n573), .B(n572), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n792), .A2(G89), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G76), .A2(n793), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT5), .B(n577), .Z(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U642 ( .A(KEYINPUT73), .B(KEYINPUT7), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n581), .B(n580), .ZN(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT74), .B(n582), .ZN(G286) );
  NAND2_X1 U646 ( .A1(G50), .A2(n796), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G62), .A2(n797), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n792), .A2(G88), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G75), .A2(n793), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT79), .B(n587), .Z(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(KEYINPUT80), .B(n590), .ZN(G166) );
  NAND2_X1 U655 ( .A1(G87), .A2(n591), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G74), .A2(G651), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U658 ( .A1(n797), .A2(n594), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n796), .A2(G49), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(G288) );
  INV_X1 U661 ( .A(G166), .ZN(G303) );
  NAND2_X1 U662 ( .A1(n793), .A2(G73), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U664 ( .A1(n792), .A2(G86), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G61), .A2(n797), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n796), .A2(G48), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT78), .B(n600), .Z(n601) );
  NOR2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n604), .A2(n603), .ZN(G305) );
  NAND2_X1 U671 ( .A1(n792), .A2(G85), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G72), .A2(n793), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U674 ( .A1(G47), .A2(n796), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G60), .A2(n797), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  OR2_X1 U677 ( .A1(n610), .A2(n609), .ZN(G290) );
  NAND2_X1 U678 ( .A1(G81), .A2(n792), .ZN(n611) );
  XOR2_X1 U679 ( .A(KEYINPUT71), .B(n611), .Z(n612) );
  XNOR2_X1 U680 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G68), .A2(n793), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n615), .B(KEYINPUT13), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G43), .A2(n796), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n797), .A2(G56), .ZN(n618) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(n618), .Z(n619) );
  NOR2_X2 U688 ( .A1(n620), .A2(n619), .ZN(n940) );
  XOR2_X1 U689 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n623) );
  NOR2_X1 U690 ( .A1(G164), .A2(G1384), .ZN(n734) );
  INV_X1 U691 ( .A(n637), .ZN(n658) );
  NAND2_X1 U692 ( .A1(n658), .A2(G1996), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G1341), .A2(n637), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT101), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n940), .A2(n627), .ZN(n642) );
  NAND2_X1 U698 ( .A1(G54), .A2(n796), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G66), .A2(n797), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n792), .A2(G92), .ZN(n631) );
  NAND2_X1 U702 ( .A1(G79), .A2(n793), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT15), .ZN(n927) );
  XNOR2_X1 U706 ( .A(n635), .B(KEYINPUT102), .ZN(n641) );
  NAND2_X1 U707 ( .A1(G1348), .A2(n677), .ZN(n639) );
  INV_X1 U708 ( .A(KEYINPUT97), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n661) );
  INV_X1 U710 ( .A(n661), .ZN(n647) );
  NAND2_X1 U711 ( .A1(G2067), .A2(n647), .ZN(n638) );
  AND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n642), .A2(n927), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n651) );
  INV_X1 U715 ( .A(G299), .ZN(n928) );
  INV_X1 U716 ( .A(G2072), .ZN(n645) );
  OR2_X1 U717 ( .A1(n661), .A2(n645), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT27), .ZN(n649) );
  INV_X1 U719 ( .A(G1956), .ZN(n1005) );
  NOR2_X1 U720 ( .A1(n647), .A2(n1005), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n928), .A2(n652), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n928), .A2(n652), .ZN(n653) );
  XOR2_X1 U725 ( .A(n653), .B(KEYINPUT28), .Z(n654) );
  NAND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n666) );
  XOR2_X1 U728 ( .A(G1961), .B(KEYINPUT95), .Z(n1000) );
  NOR2_X1 U729 ( .A1(n658), .A2(n1000), .ZN(n659) );
  XOR2_X1 U730 ( .A(KEYINPUT96), .B(n659), .Z(n664) );
  XOR2_X1 U731 ( .A(G2078), .B(KEYINPUT25), .Z(n660) );
  XNOR2_X1 U732 ( .A(KEYINPUT98), .B(n660), .ZN(n951) );
  NOR2_X1 U733 ( .A1(n951), .A2(n661), .ZN(n662) );
  XNOR2_X1 U734 ( .A(KEYINPUT99), .B(n662), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n670), .A2(G171), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n675) );
  XNOR2_X1 U738 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n669) );
  NOR2_X1 U739 ( .A1(G1966), .A2(n709), .ZN(n689) );
  NOR2_X1 U740 ( .A1(G2084), .A2(n677), .ZN(n686) );
  NAND2_X1 U741 ( .A1(n667), .A2(G8), .ZN(n668) );
  NOR2_X1 U742 ( .A1(G168), .A2(n525), .ZN(n672) );
  NOR2_X1 U743 ( .A1(G171), .A2(n670), .ZN(n671) );
  NOR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U745 ( .A(KEYINPUT31), .B(n673), .Z(n674) );
  NAND2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n690) );
  NAND2_X1 U747 ( .A1(n690), .A2(G286), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT104), .ZN(n683) );
  NOR2_X1 U749 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U750 ( .A(KEYINPUT105), .B(n678), .ZN(n681) );
  NOR2_X1 U751 ( .A1(G1971), .A2(n709), .ZN(n679) );
  NOR2_X1 U752 ( .A1(G166), .A2(n679), .ZN(n680) );
  NAND2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n684), .A2(G8), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT32), .ZN(n693) );
  NAND2_X1 U757 ( .A1(G8), .A2(n686), .ZN(n687) );
  XOR2_X1 U758 ( .A(KEYINPUT94), .B(n687), .Z(n688) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n699) );
  NOR2_X1 U762 ( .A1(G303), .A2(G1971), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n699), .A2(n695), .ZN(n936) );
  NAND2_X1 U764 ( .A1(n705), .A2(n936), .ZN(n698) );
  NAND2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n931) );
  NOR2_X1 U766 ( .A1(KEYINPUT33), .A2(n524), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n699), .A2(KEYINPUT33), .ZN(n700) );
  XOR2_X1 U768 ( .A(G1981), .B(G305), .Z(n943) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n713) );
  NOR2_X1 U770 ( .A1(G303), .A2(G2090), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n706), .A2(n709), .ZN(n711) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n707) );
  XOR2_X1 U775 ( .A(n707), .B(KEYINPUT24), .Z(n708) );
  OR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n755) );
  NAND2_X1 U779 ( .A1(G119), .A2(n885), .ZN(n715) );
  NAND2_X1 U780 ( .A1(G107), .A2(n886), .ZN(n714) );
  NAND2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U782 ( .A(KEYINPUT88), .B(n716), .Z(n722) );
  NAND2_X1 U783 ( .A1(G131), .A2(n882), .ZN(n717) );
  XOR2_X1 U784 ( .A(KEYINPUT89), .B(n717), .Z(n719) );
  NAND2_X1 U785 ( .A1(G95), .A2(n881), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U787 ( .A(KEYINPUT90), .B(n720), .Z(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n897) );
  NAND2_X1 U789 ( .A1(G1991), .A2(n897), .ZN(n723) );
  XNOR2_X1 U790 ( .A(n723), .B(KEYINPUT91), .ZN(n733) );
  NAND2_X1 U791 ( .A1(G129), .A2(n885), .ZN(n725) );
  NAND2_X1 U792 ( .A1(G117), .A2(n886), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U794 ( .A1(G105), .A2(n881), .ZN(n726) );
  XOR2_X1 U795 ( .A(KEYINPUT38), .B(n726), .Z(n727) );
  NOR2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U797 ( .A(n729), .B(KEYINPUT92), .ZN(n731) );
  NAND2_X1 U798 ( .A1(G141), .A2(n882), .ZN(n730) );
  NAND2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n894) );
  AND2_X1 U800 ( .A1(G1996), .A2(n894), .ZN(n732) );
  NOR2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n982) );
  NAND2_X1 U802 ( .A1(G160), .A2(G40), .ZN(n735) );
  NOR2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U804 ( .A(n736), .B(KEYINPUT84), .ZN(n765) );
  INV_X1 U805 ( .A(n765), .ZN(n738) );
  XOR2_X1 U806 ( .A(KEYINPUT93), .B(n738), .Z(n737) );
  NOR2_X1 U807 ( .A1(n982), .A2(n737), .ZN(n758) );
  INV_X1 U808 ( .A(n758), .ZN(n741) );
  XOR2_X1 U809 ( .A(G1986), .B(G290), .Z(n932) );
  NOR2_X1 U810 ( .A1(n932), .A2(n738), .ZN(n739) );
  XNOR2_X1 U811 ( .A(n739), .B(KEYINPUT85), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n753) );
  XNOR2_X1 U813 ( .A(G2067), .B(KEYINPUT37), .ZN(n763) );
  NAND2_X1 U814 ( .A1(G104), .A2(n881), .ZN(n743) );
  NAND2_X1 U815 ( .A1(G140), .A2(n882), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U817 ( .A(KEYINPUT34), .B(n744), .ZN(n751) );
  NAND2_X1 U818 ( .A1(n885), .A2(G128), .ZN(n745) );
  XNOR2_X1 U819 ( .A(n745), .B(KEYINPUT86), .ZN(n747) );
  NAND2_X1 U820 ( .A1(G116), .A2(n886), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U822 ( .A(KEYINPUT87), .B(n748), .ZN(n749) );
  XNOR2_X1 U823 ( .A(KEYINPUT35), .B(n749), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U825 ( .A(KEYINPUT36), .B(n752), .ZN(n865) );
  NOR2_X1 U826 ( .A1(n763), .A2(n865), .ZN(n981) );
  OR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n768) );
  NOR2_X1 U828 ( .A1(G1996), .A2(n894), .ZN(n988) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n756) );
  NOR2_X1 U830 ( .A1(G1991), .A2(n897), .ZN(n978) );
  NOR2_X1 U831 ( .A1(n756), .A2(n978), .ZN(n757) );
  NOR2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n988), .A2(n759), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT39), .ZN(n762) );
  INV_X1 U835 ( .A(n981), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U837 ( .A1(n763), .A2(n865), .ZN(n985) );
  NAND2_X1 U838 ( .A1(n764), .A2(n985), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n769), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U843 ( .A(KEYINPUT18), .B(KEYINPUT76), .Z(n771) );
  NAND2_X1 U844 ( .A1(G123), .A2(n885), .ZN(n770) );
  XNOR2_X1 U845 ( .A(n771), .B(n770), .ZN(n775) );
  NAND2_X1 U846 ( .A1(n886), .A2(G111), .ZN(n773) );
  NAND2_X1 U847 ( .A1(G99), .A2(n881), .ZN(n772) );
  NAND2_X1 U848 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U849 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U850 ( .A1(G135), .A2(n882), .ZN(n776) );
  NAND2_X1 U851 ( .A1(n777), .A2(n776), .ZN(n975) );
  XNOR2_X1 U852 ( .A(G2096), .B(n975), .ZN(n778) );
  OR2_X1 U853 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  INV_X1 U856 ( .A(G82), .ZN(G220) );
  NAND2_X1 U857 ( .A1(G7), .A2(G661), .ZN(n779) );
  XNOR2_X1 U858 ( .A(n779), .B(KEYINPUT70), .ZN(n780) );
  XNOR2_X1 U859 ( .A(KEYINPUT10), .B(n780), .ZN(G223) );
  INV_X1 U860 ( .A(G223), .ZN(n832) );
  NAND2_X1 U861 ( .A1(n832), .A2(G567), .ZN(n781) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  NAND2_X1 U863 ( .A1(n940), .A2(G860), .ZN(G153) );
  INV_X1 U864 ( .A(G171), .ZN(G301) );
  NAND2_X1 U865 ( .A1(G868), .A2(G301), .ZN(n783) );
  INV_X1 U866 ( .A(G868), .ZN(n817) );
  NAND2_X1 U867 ( .A1(n927), .A2(n817), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(G284) );
  NAND2_X1 U869 ( .A1(G868), .A2(G286), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G299), .A2(n817), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(G297) );
  INV_X1 U872 ( .A(G860), .ZN(n804) );
  NAND2_X1 U873 ( .A1(n804), .A2(G559), .ZN(n786) );
  INV_X1 U874 ( .A(n927), .ZN(n802) );
  NAND2_X1 U875 ( .A1(n786), .A2(n802), .ZN(n787) );
  XNOR2_X1 U876 ( .A(n787), .B(KEYINPUT75), .ZN(n788) );
  XOR2_X1 U877 ( .A(KEYINPUT16), .B(n788), .Z(G148) );
  NAND2_X1 U878 ( .A1(n802), .A2(G868), .ZN(n789) );
  NOR2_X1 U879 ( .A1(G559), .A2(n789), .ZN(n791) );
  AND2_X1 U880 ( .A1(n817), .A2(n940), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U882 ( .A1(n792), .A2(G93), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G80), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G55), .A2(n796), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G67), .A2(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n816) );
  NAND2_X1 U889 ( .A1(G559), .A2(n802), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n803), .B(n940), .ZN(n814) );
  NAND2_X1 U891 ( .A1(n804), .A2(n814), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n805), .B(KEYINPUT77), .ZN(n806) );
  XOR2_X1 U893 ( .A(n816), .B(n806), .Z(G145) );
  XNOR2_X1 U894 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n808) );
  XNOR2_X1 U895 ( .A(G288), .B(KEYINPUT81), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n809) );
  XOR2_X1 U897 ( .A(n816), .B(n809), .Z(n811) );
  XNOR2_X1 U898 ( .A(G290), .B(n928), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(G166), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n813), .B(G305), .ZN(n900) );
  XNOR2_X1 U902 ( .A(n814), .B(n900), .ZN(n815) );
  NAND2_X1 U903 ( .A1(n815), .A2(G868), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n821), .ZN(n822) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n823), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n824) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n824), .Z(n825) );
  NOR2_X1 U914 ( .A1(G218), .A2(n825), .ZN(n826) );
  NAND2_X1 U915 ( .A1(G96), .A2(n826), .ZN(n922) );
  NAND2_X1 U916 ( .A1(n922), .A2(G2106), .ZN(n830) );
  NAND2_X1 U917 ( .A1(G69), .A2(G120), .ZN(n827) );
  NOR2_X1 U918 ( .A1(G237), .A2(n827), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G108), .A2(n828), .ZN(n923) );
  NAND2_X1 U920 ( .A1(n923), .A2(G567), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n830), .A2(n829), .ZN(n837) );
  NAND2_X1 U922 ( .A1(G483), .A2(G661), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n837), .A2(n831), .ZN(n836) );
  NAND2_X1 U924 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XOR2_X1 U926 ( .A(KEYINPUT109), .B(n833), .Z(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U928 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U931 ( .A(n837), .ZN(G319) );
  XNOR2_X1 U932 ( .A(G1996), .B(G2474), .ZN(n847) );
  XOR2_X1 U933 ( .A(G1981), .B(G1961), .Z(n839) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1966), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1956), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U940 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(G229) );
  XOR2_X1 U943 ( .A(G2100), .B(G2096), .Z(n849) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2072), .Z(n851) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U949 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U952 ( .A1(n885), .A2(G124), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U954 ( .A1(G136), .A2(n882), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n859), .B(KEYINPUT111), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G100), .A2(n881), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U959 ( .A1(n886), .A2(G112), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT112), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G162), .B(n865), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n866), .B(n975), .ZN(n870) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n868) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(n870), .B(n869), .Z(n880) );
  NAND2_X1 U968 ( .A1(G130), .A2(n885), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G118), .A2(n886), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G106), .A2(n881), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G142), .A2(n882), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n875), .Z(n876) );
  NOR2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U976 ( .A(G160), .B(n878), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n893) );
  NAND2_X1 U978 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U981 ( .A1(G127), .A2(n885), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G115), .A2(n886), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U986 ( .A(KEYINPUT113), .B(n892), .Z(n971) );
  XOR2_X1 U987 ( .A(n893), .B(n971), .Z(n896) );
  XOR2_X1 U988 ( .A(n894), .B(G164), .Z(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U991 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G286), .B(n900), .ZN(n902) );
  XNOR2_X1 U993 ( .A(G171), .B(n940), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U995 ( .A(n927), .B(KEYINPUT116), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G37), .A2(n905), .ZN(G397) );
  XNOR2_X1 U998 ( .A(G2451), .B(G2446), .ZN(n915) );
  XOR2_X1 U999 ( .A(G2430), .B(KEYINPUT108), .Z(n907) );
  XNOR2_X1 U1000 ( .A(G2454), .B(G2435), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1002 ( .A(G2438), .B(KEYINPUT107), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G2443), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1009 ( .A1(n916), .A2(G14), .ZN(n924) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n924), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(G225) );
  XNOR2_X1 U1016 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G120), .ZN(G236) );
  INV_X1 U1019 ( .A(G96), .ZN(G221) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(G325) );
  INV_X1 U1022 ( .A(G325), .ZN(G261) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  INV_X1 U1024 ( .A(n924), .ZN(G401) );
  XNOR2_X1 U1025 ( .A(G1961), .B(G171), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n938) );
  XOR2_X1 U1028 ( .A(n927), .B(G1348), .Z(n930) );
  XNOR2_X1 U1029 ( .A(n928), .B(G1956), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(n939), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n940), .B(G1341), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G168), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1040 ( .A(KEYINPUT57), .B(n945), .Z(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n949) );
  XOR2_X1 U1042 ( .A(G16), .B(KEYINPUT56), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(KEYINPUT125), .B(n950), .ZN(n970) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n963) );
  XNOR2_X1 U1046 ( .A(n951), .B(G27), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G32), .B(G1996), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(n954), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G1991), .B(G25), .Z(n959) );
  NAND2_X1 U1055 ( .A1(G28), .A2(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n963), .B(n962), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G2084), .B(G34), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT54), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G35), .B(G2090), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n1026) );
  INV_X1 U1063 ( .A(KEYINPUT55), .ZN(n998) );
  OR2_X1 U1064 ( .A1(n1026), .A2(n998), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n1033) );
  XOR2_X1 U1066 ( .A(G2072), .B(n971), .Z(n973) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT50), .B(n974), .ZN(n995) );
  XNOR2_X1 U1070 ( .A(G160), .B(G2084), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(KEYINPUT118), .B(n979), .Z(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n984), .B(KEYINPUT119), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n993) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1080 ( .A(KEYINPUT51), .B(n989), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(n991), .B(n990), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT52), .B(n996), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n999), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G21), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(n1000), .B(G5), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1014) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(G4), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1004), .B(n1003), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(G20), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT60), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1022) );
  XNOR2_X1 U1102 ( .A(G1986), .B(G24), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT127), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1023), .Z(n1024) );
  NOR2_X1 U1111 ( .A1(G16), .A2(n1024), .ZN(n1029) );
  NOR2_X1 U1112 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(G11), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(n1034), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

