//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n212), .B1(new_n201), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G244), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n214), .B1(G77), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G97), .A2(G257), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n211), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NOR4_X1   g0034(.A1(new_n224), .A2(new_n226), .A3(new_n229), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n204), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n232), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n252), .B1(new_n253), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n233), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n258), .A2(new_n260), .B1(new_n201), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT68), .A2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT68), .A2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI211_X1 g0078(.A(G1), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n233), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n213), .ZN(new_n286));
  OR3_X1    g0086(.A1(new_n279), .A2(new_n286), .A3(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n288), .B2(new_n290), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n281), .A2(new_n282), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n233), .ZN(new_n298));
  MUX2_X1   g0098(.A(G222), .B(G223), .S(G1698), .Z(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n298), .C1(new_n294), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT69), .B1(new_n279), .B2(new_n286), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n287), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n271), .B(new_n272), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(G200), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n311), .A3(new_n307), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n312), .A2(KEYINPUT74), .A3(KEYINPUT10), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT74), .B1(new_n312), .B2(KEYINPUT10), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n289), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n281), .A2(KEYINPUT3), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT70), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n213), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n321), .B(new_n323), .C1(G232), .C2(new_n322), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n283), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n279), .ZN(new_n327));
  INV_X1    g0127(.A(G238), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n285), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n316), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n326), .A2(KEYINPUT13), .A3(new_n279), .A4(new_n329), .ZN(new_n332));
  OAI21_X1  g0132(.A(G169), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n331), .A2(new_n332), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(G169), .C1(new_n331), .C2(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n255), .A2(new_n201), .B1(new_n232), .B2(G68), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n256), .A2(new_n295), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n260), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT11), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n263), .A2(new_n203), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT12), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n259), .A2(new_n233), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(KEYINPUT72), .A3(new_n262), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n263), .B2(new_n260), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n266), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G68), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n343), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G200), .B1(new_n331), .B2(new_n332), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n335), .A2(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n302), .A2(G179), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n302), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n269), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n315), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n257), .A2(new_n262), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n267), .B2(new_n257), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n230), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G20), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT75), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n254), .A2(G159), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(KEYINPUT75), .A3(G20), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT3), .B(G33), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n376), .A2(new_n377), .A3(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n319), .A2(new_n232), .A3(new_n320), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n380), .B2(new_n203), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n377), .B1(new_n376), .B2(G20), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n288), .A2(new_n290), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n203), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n346), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n367), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n213), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n376), .B(new_n393), .C1(G223), .C2(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n298), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n285), .A2(new_n237), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n277), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n261), .B(G274), .C1(new_n400), .C2(G45), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n283), .B1(new_n394), .B2(new_n395), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n404), .A2(new_n279), .A3(new_n398), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G179), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n392), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(new_n407), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n391), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n397), .A2(new_n399), .A3(new_n303), .A4(new_n401), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n405), .B2(G200), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n294), .B2(new_n232), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n415), .B2(new_n378), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT16), .B1(new_n416), .B2(new_n375), .ZN(new_n417));
  INV_X1    g0217(.A(new_n388), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n375), .A2(new_n418), .A3(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n260), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n366), .B(new_n414), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT76), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n391), .A2(KEYINPUT76), .A3(new_n414), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n391), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT17), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n421), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n412), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n257), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(KEYINPUT71), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(KEYINPUT71), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT15), .B(G87), .Z(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n433), .B(new_n434), .C1(new_n436), .C2(new_n256), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n260), .B1(G77), .B2(new_n350), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n263), .A2(new_n295), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n328), .A2(G1698), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G232), .B2(G1698), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n283), .B1(new_n321), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G107), .B2(new_n321), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n283), .A2(new_n215), .A3(new_n284), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n401), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n361), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(G179), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n446), .A2(new_n303), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(G200), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n439), .A3(new_n438), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n430), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n364), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n220), .A2(G1698), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n288), .A3(new_n290), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT90), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n376), .A2(G257), .A3(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n455), .A2(new_n288), .A3(new_n290), .A4(KEYINPUT90), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n298), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n261), .A2(G45), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(KEYINPUT5), .B2(new_n282), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n275), .A2(new_n466), .A3(new_n276), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n467), .A3(G274), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n298), .B1(new_n465), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G264), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n463), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT91), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n462), .A2(new_n298), .B1(new_n469), .B2(G264), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT91), .A3(new_n468), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n303), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G200), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n219), .A2(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT22), .B1(new_n321), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G116), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G20), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n232), .A2(KEYINPUT22), .A3(G87), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n376), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT87), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n490), .A2(new_n486), .A3(new_n487), .A4(G20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT23), .B1(new_n232), .B2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n485), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT88), .B1(new_n481), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n480), .B1(new_n292), .B2(new_n293), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT22), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n485), .A2(new_n492), .A3(new_n493), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT88), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n501), .A3(KEYINPUT24), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT24), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT88), .B(new_n503), .C1(new_n481), .C2(new_n494), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n260), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n263), .A2(new_n260), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n281), .A2(G1), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(new_n487), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n262), .A2(G107), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT89), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT25), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n479), .A2(new_n505), .A3(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n502), .A2(new_n260), .A3(new_n504), .ZN(new_n518));
  INV_X1    g0318(.A(new_n516), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n361), .B1(new_n473), .B2(new_n475), .ZN(new_n520));
  INV_X1    g0320(.A(G179), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n471), .A2(new_n521), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n288), .A2(new_n290), .A3(G244), .A4(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n376), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n376), .A2(G238), .A3(new_n322), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n482), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n298), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(new_n464), .C1(new_n297), .C2(new_n233), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n273), .B2(new_n464), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(KEYINPUT81), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n361), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT81), .B1(new_n530), .B2(new_n533), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n535), .B(new_n532), .C1(new_n529), .C2(new_n298), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n521), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n232), .B1(new_n325), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n207), .A2(G87), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n376), .A2(new_n232), .A3(G68), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n256), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(KEYINPUT19), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n260), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n435), .A2(new_n262), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(new_n509), .C2(new_n436), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n538), .A2(new_n541), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n536), .A2(G200), .A3(new_n537), .ZN(new_n557));
  OAI21_X1  g0357(.A(G190), .B1(new_n539), .B2(new_n540), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n506), .A2(G87), .A3(new_n508), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n552), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n517), .A2(new_n523), .A3(new_n556), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n276), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n563), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n278), .A2(G1), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n466), .B2(G41), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n283), .B(G257), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n468), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n570), .A3(new_n468), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(G250), .B1(new_n292), .B2(new_n293), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n322), .B1(new_n573), .B2(KEYINPUT4), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT4), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G1698), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(new_n576), .C1(new_n292), .C2(new_n293), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT4), .B1(new_n376), .B2(G244), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G283), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n574), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n521), .B(new_n572), .C1(new_n583), .C2(new_n283), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n574), .A2(new_n582), .ZN(new_n586));
  INV_X1    g0386(.A(G244), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n319), .B2(new_n320), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n578), .B1(new_n588), .B2(new_n576), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n283), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n361), .B1(new_n590), .B2(new_n568), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n262), .A2(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n254), .A2(G77), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n549), .A2(new_n487), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(new_n206), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n596), .B2(KEYINPUT6), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G20), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n593), .B(new_n598), .C1(new_n380), .C2(new_n487), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n599), .B2(new_n260), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n509), .A2(new_n549), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n220), .B1(new_n319), .B2(new_n320), .ZN(new_n604));
  OAI21_X1  g0404(.A(G1698), .B1(new_n604), .B2(new_n575), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n589), .A3(new_n581), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n298), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT79), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n521), .A4(new_n572), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n585), .A2(new_n591), .A3(new_n603), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n572), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G200), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n568), .B1(new_n606), .B2(new_n298), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G190), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n600), .A3(new_n602), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  INV_X1    g0417(.A(G116), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n618), .B(new_n507), .C1(new_n347), .C2(new_n349), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n259), .A2(new_n233), .B1(G20), .B2(new_n618), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n581), .B(new_n232), .C1(G33), .C2(new_n549), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT20), .B1(new_n620), .B2(new_n621), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(G116), .B2(new_n262), .ZN(new_n624));
  OAI21_X1  g0424(.A(G169), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n283), .B(G270), .C1(new_n564), .C2(new_n566), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n468), .ZN(new_n627));
  XOR2_X1   g0427(.A(KEYINPUT84), .B(G303), .Z(new_n628));
  NAND3_X1  g0428(.A1(new_n319), .A2(new_n320), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT83), .ZN(new_n630));
  NAND2_X1  g0430(.A1(G264), .A2(G1698), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n386), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n376), .A2(KEYINPUT83), .A3(G264), .A4(G1698), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n376), .A2(G257), .A3(new_n322), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n627), .B1(new_n635), .B2(new_n298), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n617), .B1(new_n625), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT86), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT86), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(new_n617), .C1(new_n625), .C2(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(G190), .ZN(new_n642));
  INV_X1    g0442(.A(new_n623), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n620), .A2(KEYINPUT20), .A3(new_n621), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n643), .A2(new_n644), .B1(new_n618), .B2(new_n263), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n347), .A2(new_n349), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(G116), .A3(new_n508), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n642), .B(new_n649), .C1(new_n477), .C2(new_n636), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n635), .A2(new_n298), .ZN(new_n651));
  INV_X1    g0451(.A(new_n627), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(KEYINPUT21), .A3(G169), .A4(new_n648), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n636), .A2(new_n648), .A3(G179), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n654), .A2(KEYINPUT85), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT85), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n641), .B(new_n650), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n562), .A2(new_n616), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n454), .A2(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n363), .ZN(new_n661));
  INV_X1    g0461(.A(new_n412), .ZN(new_n662));
  INV_X1    g0462(.A(new_n449), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n358), .A2(new_n663), .B1(new_n339), .B2(new_n352), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n428), .B1(new_n426), .B2(KEYINPUT17), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n661), .B1(new_n666), .B2(new_n315), .ZN(new_n667));
  INV_X1    g0467(.A(new_n454), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT92), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n654), .A2(new_n655), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n641), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n475), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT91), .B1(new_n474), .B2(new_n468), .ZN(new_n673));
  OAI21_X1  g0473(.A(G169), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n522), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n505), .B2(new_n516), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n669), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n641), .A4(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n534), .A2(new_n361), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n541), .A2(new_n555), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n534), .A2(G200), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n558), .A2(new_n560), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n610), .A3(new_n615), .A4(new_n517), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n609), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n606), .A2(new_n298), .B1(new_n569), .B2(new_n571), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n608), .B1(new_n688), .B2(new_n521), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n591), .A2(new_n603), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n684), .A2(new_n690), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n556), .A2(new_n561), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n610), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n695), .A3(new_n681), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n693), .A2(new_n695), .A3(KEYINPUT93), .A4(new_n681), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n686), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n667), .B1(new_n668), .B2(new_n700), .ZN(G369));
  INV_X1    g0501(.A(G13), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G20), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n261), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G213), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n649), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n671), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n658), .A2(KEYINPUT94), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n658), .A2(KEYINPUT94), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n712), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n505), .A2(new_n516), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n709), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n517), .A2(new_n523), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n676), .A2(new_n709), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT95), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n716), .A2(new_n722), .A3(G330), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n641), .B1(new_n656), .B2(new_n657), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n710), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n719), .B2(new_n720), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n523), .A2(new_n709), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n723), .A2(new_n730), .A3(new_n732), .ZN(G399));
  INV_X1    g0533(.A(new_n227), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n400), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n546), .A2(new_n618), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(G1), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n231), .B2(new_n736), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n536), .A2(new_n537), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n636), .A2(G179), .A3(new_n474), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(new_n743), .A3(new_n613), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT96), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(G179), .B1(new_n530), .B2(new_n533), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n611), .A2(new_n471), .A3(new_n653), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n744), .B2(new_n746), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(new_n746), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n710), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n717), .B1(new_n476), .B2(new_n478), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n755), .A2(new_n694), .A3(new_n676), .ZN(new_n756));
  INV_X1    g0556(.A(new_n616), .ZN(new_n757));
  INV_X1    g0557(.A(new_n658), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n756), .A2(new_n757), .A3(new_n758), .A4(new_n710), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n754), .B1(new_n759), .B2(KEYINPUT31), .ZN(new_n760));
  INV_X1    g0560(.A(new_n752), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(new_n750), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G330), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT29), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n700), .B2(new_n709), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n681), .A2(new_n683), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT26), .B1(new_n610), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n690), .A2(new_n692), .A3(new_n556), .A4(new_n561), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n681), .B(new_n771), .C1(new_n772), .C2(KEYINPUT26), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n724), .A2(new_n676), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n685), .ZN(new_n775));
  OAI211_X1 g0575(.A(KEYINPUT29), .B(new_n710), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n767), .B1(new_n769), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n741), .B1(new_n777), .B2(G1), .ZN(G364));
  NAND2_X1  g0578(.A1(new_n703), .A2(G45), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n736), .A2(G1), .A3(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n233), .B1(G20), .B2(new_n361), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n232), .A2(G190), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(new_n521), .A3(new_n477), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT101), .B(G159), .Z(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n477), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n792), .A2(KEYINPUT32), .B1(new_n487), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n303), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(G50), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n232), .A2(new_n303), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n521), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G58), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n303), .A2(G179), .A3(G200), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n232), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n805), .A2(KEYINPUT102), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(KEYINPUT102), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n792), .A2(KEYINPUT32), .B1(new_n809), .B2(G97), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n799), .A2(new_n793), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G87), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n796), .A2(G190), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n203), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n800), .A2(new_n784), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n294), .B(new_n816), .C1(G77), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n798), .A2(new_n803), .A3(new_n810), .A4(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G329), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n788), .A2(new_n823), .B1(new_n824), .B2(new_n794), .ZN(new_n825));
  INV_X1    g0625(.A(new_n805), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n822), .B(new_n825), .C1(G294), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n802), .A2(G322), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n797), .A2(G326), .ZN(new_n829));
  INV_X1    g0629(.A(G303), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n811), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n831), .B(new_n321), .C1(new_n814), .C2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n783), .B1(new_n820), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(G13), .A2(G33), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT98), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n232), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n782), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n734), .A2(new_n376), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n250), .B2(new_n278), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n231), .A2(G45), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(G116), .B2(new_n227), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n294), .A2(new_n734), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G355), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT97), .Z(new_n848));
  AOI21_X1  g0648(.A(new_n835), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n781), .B(new_n849), .C1(new_n716), .C2(new_n839), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n716), .B(G330), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n781), .ZN(G396));
  OR2_X1    g0652(.A1(new_n679), .A2(new_n685), .ZN(new_n853));
  INV_X1    g0653(.A(new_n681), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n772), .B2(KEYINPUT26), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT93), .B1(new_n855), .B2(new_n693), .ZN(new_n856));
  INV_X1    g0656(.A(new_n699), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n440), .A2(new_n709), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n449), .A2(new_n452), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT104), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT104), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n449), .A2(new_n859), .A3(new_n862), .A4(new_n452), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(new_n710), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n663), .A2(new_n709), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n700), .B2(new_n709), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n767), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n874), .B(new_n780), .C1(new_n767), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n869), .A2(new_n837), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n814), .A2(G150), .B1(new_n797), .B2(G137), .ZN(new_n877));
  INV_X1    g0677(.A(G143), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n877), .B1(new_n878), .B2(new_n801), .C1(new_n817), .C2(new_n790), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT34), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n794), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n880), .B1(G68), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n826), .A2(G58), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n376), .B1(new_n811), .B2(new_n201), .ZN(new_n885));
  INV_X1    g0685(.A(new_n788), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(G132), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n794), .A2(new_n219), .ZN(new_n889));
  INV_X1    g0689(.A(new_n797), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n890), .A2(new_n830), .B1(new_n817), .B2(new_n618), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(G283), .B2(new_n814), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT103), .Z(new_n893));
  AOI211_X1 g0693(.A(new_n889), .B(new_n893), .C1(G294), .C2(new_n802), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n549), .B2(new_n808), .C1(new_n821), .C2(new_n788), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n294), .B1(new_n487), .B2(new_n811), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n782), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n837), .A2(new_n782), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n295), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n876), .A2(new_n781), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n875), .A2(new_n901), .ZN(G384));
  NAND2_X1  g0702(.A1(new_n352), .A2(new_n709), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n353), .A2(new_n358), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n339), .A2(new_n352), .A3(new_n709), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n747), .A2(new_n750), .ZN(new_n907));
  INV_X1    g0707(.A(new_n753), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT31), .B(new_n709), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n868), .B(new_n906), .C1(new_n760), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n423), .A2(new_n424), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n391), .A2(new_n707), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n391), .A2(new_n410), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n410), .A2(new_n707), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n389), .B1(new_n920), .B2(KEYINPUT16), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT106), .B(new_n382), .C1(new_n384), .C2(new_n388), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n260), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n366), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n423), .A2(new_n424), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n917), .A2(new_n918), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  INV_X1    g0726(.A(new_n707), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n926), .B1(new_n430), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT38), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(KEYINPUT107), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT107), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n927), .B(new_n924), .C1(new_n665), .C2(new_n412), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT38), .A3(new_n926), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n912), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n934), .A2(KEYINPUT38), .A3(new_n926), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n915), .B1(new_n665), .B2(new_n412), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n421), .B1(new_n391), .B2(new_n410), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT37), .B1(new_n942), .B2(new_n915), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n917), .B2(new_n918), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT40), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n911), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(G330), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT31), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n659), .B2(new_n710), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n909), .B1(new_n951), .B2(new_n754), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n454), .A2(G330), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n947), .B1(new_n937), .B2(new_n938), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n454), .A2(new_n952), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n949), .A2(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n931), .ZN(new_n957));
  XOR2_X1   g0757(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n958));
  AND2_X1   g0758(.A1(new_n941), .A2(new_n944), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n935), .B(new_n958), .C1(new_n959), .C2(KEYINPUT38), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n353), .A2(new_n709), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n906), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n449), .A2(new_n709), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n866), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n931), .A3(new_n936), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n662), .A2(new_n927), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n956), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n769), .A2(new_n454), .A3(new_n776), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n667), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n261), .B2(new_n703), .ZN(new_n976));
  OAI211_X1 g0776(.A(G20), .B(new_n280), .C1(new_n597), .C2(KEYINPUT35), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n618), .B(new_n977), .C1(KEYINPUT35), .C2(new_n597), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT36), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n368), .A2(G77), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n231), .A2(new_n980), .B1(G50), .B2(new_n203), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(G1), .A3(new_n702), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n976), .A2(new_n979), .A3(new_n982), .ZN(G367));
  NAND2_X1  g0783(.A1(new_n730), .A2(new_n732), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n603), .A2(new_n709), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n615), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n610), .ZN(new_n987));
  INV_X1    g0787(.A(new_n610), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n710), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n984), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n722), .A2(new_n726), .A3(new_n987), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n995), .A3(new_n989), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n560), .A2(new_n710), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT109), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(new_n770), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n854), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n996), .A2(KEYINPUT43), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n996), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n723), .A2(new_n990), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n735), .B(KEYINPUT41), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n716), .A2(new_n722), .A3(G330), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n722), .B1(new_n716), .B2(G330), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n725), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n716), .A2(G330), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n722), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n723), .A3(new_n726), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n769), .A2(new_n776), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n763), .B1(new_n951), .B2(new_n754), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(G330), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT110), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT110), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n777), .A2(new_n1025), .A3(new_n1018), .A4(new_n1014), .ZN(new_n1026));
  AOI21_X1  g0826(.A(KEYINPUT44), .B1(new_n984), .B2(new_n990), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1028), .B(new_n991), .C1(new_n730), .C2(new_n732), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n730), .A2(new_n732), .A3(new_n991), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT45), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n723), .B1(new_n1027), .B2(new_n1029), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1033), .A2(new_n1032), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n1012), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1024), .A2(new_n1026), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1011), .B1(new_n1037), .B2(new_n777), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n779), .A2(G1), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT111), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1009), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n788), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1044), .A2(KEYINPUT112), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n817), .A2(new_n824), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT46), .B1(new_n812), .B2(G116), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(G294), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n805), .A2(new_n487), .B1(new_n815), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n628), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n386), .B1(new_n794), .B2(new_n549), .C1(new_n1051), .C2(new_n801), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(KEYINPUT112), .C2(new_n1044), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1048), .B(new_n1053), .C1(new_n821), .C2(new_n890), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n818), .A2(G50), .B1(new_n789), .B2(new_n814), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n809), .A2(G68), .B1(KEYINPUT113), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n886), .A2(G137), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n294), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n794), .A2(new_n295), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n890), .A2(new_n878), .B1(new_n801), .B2(new_n253), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G58), .C2(new_n812), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1054), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT114), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT47), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n782), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n999), .A2(new_n840), .A3(new_n1000), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n842), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n841), .B1(new_n227), .B2(new_n436), .C1(new_n243), .C2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n781), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1041), .A2(KEYINPUT115), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT115), .B1(new_n1041), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(G387));
  AOI21_X1  g0876(.A(new_n780), .B1(new_n1016), .B2(new_n840), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n240), .A2(new_n278), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(new_n842), .B1(new_n737), .B2(new_n846), .ZN(new_n1079));
  AOI21_X1  g0879(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n431), .A2(new_n201), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n738), .B(new_n1080), .C1(new_n1081), .C2(KEYINPUT50), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(KEYINPUT50), .B2(new_n1081), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1079), .A2(new_n1083), .B1(G107), .B2(new_n227), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n841), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n814), .A2(G311), .B1(new_n797), .B2(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n1042), .B2(new_n801), .C1(new_n1051), .C2(new_n817), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT48), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n805), .A2(new_n824), .B1(new_n811), .B2(new_n1049), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT118), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT49), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n886), .A2(G326), .B1(G116), .B2(new_n882), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n386), .A3(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n808), .A2(new_n436), .B1(new_n201), .B2(new_n801), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT116), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n882), .A2(G97), .B1(G159), .B2(new_n797), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n812), .A2(G77), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n818), .A2(G68), .B1(new_n431), .B2(new_n814), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n376), .B1(new_n788), .B2(new_n253), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n782), .B1(new_n1096), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1077), .A2(new_n1085), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1040), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n735), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1107), .B1(new_n1019), .B2(new_n1108), .C1(new_n1110), .C2(new_n1111), .ZN(G393));
  AND2_X1   g0912(.A1(new_n1036), .A2(new_n1034), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1037), .B(new_n735), .C1(new_n1113), .C2(new_n1111), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n841), .B1(new_n549), .B2(new_n227), .C1(new_n247), .C2(new_n1069), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n889), .B1(G68), .B2(new_n812), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n201), .B2(new_n815), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n386), .B(new_n1117), .C1(new_n431), .C2(new_n818), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n808), .A2(new_n295), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G143), .B2(new_n886), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n802), .A2(G159), .B1(G150), .B2(new_n797), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT51), .Z(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n802), .A2(G311), .B1(G317), .B2(new_n797), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT52), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G283), .B2(new_n812), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n818), .A2(G294), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n886), .A2(G322), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1051), .A2(new_n815), .B1(new_n487), .B2(new_n794), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n321), .B(new_n1129), .C1(G116), .C2(new_n826), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n783), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n780), .B(new_n1132), .C1(new_n990), .C2(new_n840), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1113), .A2(new_n1040), .B1(new_n1115), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1114), .A2(new_n1134), .ZN(G390));
  AND2_X1   g0935(.A1(new_n957), .A2(new_n960), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n837), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n812), .A2(G150), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1138), .A2(KEYINPUT53), .ZN(new_n1139));
  INV_X1    g0939(.A(G125), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n788), .A2(new_n1140), .B1(KEYINPUT53), .B2(new_n1138), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  AOI211_X1 g0942(.A(new_n1139), .B(new_n1141), .C1(new_n818), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n814), .A2(G137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n809), .A2(G159), .ZN(new_n1145));
  INV_X1    g0945(.A(G132), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n801), .A2(new_n1146), .B1(new_n794), .B2(new_n201), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n294), .B(new_n1147), .C1(G128), .C2(new_n797), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n788), .A2(new_n1049), .B1(new_n203), .B2(new_n794), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT121), .Z(new_n1151));
  OAI22_X1  g0951(.A1(new_n890), .A2(new_n824), .B1(new_n817), .B2(new_n549), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G107), .B2(new_n814), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT120), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n321), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n802), .A2(G116), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1151), .A2(new_n1155), .A3(new_n813), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1149), .B1(new_n1157), .B2(new_n1119), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n782), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n899), .A2(new_n257), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1137), .A2(new_n781), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1021), .A2(G330), .A3(new_n868), .A4(new_n906), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n865), .B(new_n710), .C1(new_n773), .C2(new_n775), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n964), .B1(new_n1163), .B2(new_n966), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n962), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n940), .B2(new_n945), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n866), .A2(new_n966), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n962), .B1(new_n1169), .B2(new_n906), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1162), .B(new_n1168), .C1(new_n1170), .C2(new_n961), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n698), .A2(new_n699), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n709), .B1(new_n1172), .B2(new_n853), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n965), .B1(new_n1173), .B2(new_n865), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1165), .B1(new_n1174), .B2(new_n964), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1167), .B1(new_n1136), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n952), .A2(G330), .A3(new_n868), .A4(new_n906), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1161), .B1(new_n1178), .B2(new_n1108), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1171), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n957), .B(new_n960), .C1(new_n967), .C2(new_n962), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n1181), .B2(new_n1168), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n868), .C1(new_n760), .C2(new_n910), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n964), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1163), .A2(new_n966), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1185), .A2(new_n1162), .A3(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G330), .B(new_n868), .C1(new_n760), .C2(new_n764), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n964), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1189), .A2(new_n1177), .B1(new_n866), .B2(new_n966), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n973), .A2(new_n953), .A3(new_n667), .ZN(new_n1192));
  OAI21_X1  g0992(.A(KEYINPUT119), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(new_n1162), .A3(new_n1186), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n912), .A2(G330), .B1(new_n964), .B2(new_n1188), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n1174), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT119), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n973), .A2(new_n953), .A3(new_n667), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1193), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n736), .B1(new_n1183), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1178), .A2(new_n1199), .A3(new_n1193), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1179), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(G378));
  NAND2_X1  g1004(.A1(new_n269), .A2(new_n927), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n315), .A2(new_n363), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n315), .B2(new_n363), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OR3_X1    g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n837), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n400), .A2(new_n376), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n549), .B2(new_n815), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n809), .A2(G68), .B1(G107), .B2(new_n802), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n618), .B2(new_n890), .C1(new_n436), .C2(new_n817), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G283), .B2(new_n886), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n202), .B2(new_n794), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1216), .B(new_n1220), .C1(G77), .C2(new_n812), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G128), .A2(new_n802), .B1(new_n818), .B2(G137), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n812), .A2(new_n1142), .B1(G132), .B2(new_n814), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1140), .C2(new_n890), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G150), .B2(new_n809), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n882), .A2(new_n789), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G33), .A2(G41), .ZN(new_n1230));
  XOR2_X1   g1030(.A(KEYINPUT122), .B(G124), .Z(new_n1231));
  NAND2_X1  g1031(.A1(new_n886), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n1215), .A2(G50), .A3(new_n1230), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1222), .A2(new_n1223), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n782), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n899), .A2(new_n201), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n781), .A2(new_n1214), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n954), .A2(G330), .A3(new_n1212), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1212), .B1(new_n954), .B2(G330), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n971), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n963), .A2(new_n968), .A3(new_n970), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n949), .A2(new_n1213), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n954), .A2(G330), .A3(new_n1212), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1238), .B1(new_n1246), .B2(new_n1040), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1181), .A2(new_n1168), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1177), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1197), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1171), .B(new_n1250), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1253), .A2(new_n1198), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n735), .B1(new_n1254), .B2(KEYINPUT57), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1178), .B1(new_n1199), .B2(new_n1193), .ZN(new_n1256));
  OAI211_X1 g1056(.A(KEYINPUT57), .B(new_n1246), .C1(new_n1256), .C2(new_n1192), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1247), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1259), .B(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(G375));
  NAND2_X1  g1062(.A1(new_n1196), .A2(new_n1040), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n817), .A2(new_n487), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n321), .B1(new_n886), .B2(G303), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n618), .B2(new_n815), .C1(new_n1049), .C2(new_n890), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(new_n1266), .C1(G283), .C2(new_n802), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1060), .B1(new_n809), .B2(new_n435), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(new_n549), .C2(new_n811), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT125), .Z(new_n1270));
  AOI22_X1  g1070(.A1(new_n809), .A2(G50), .B1(G150), .B2(new_n818), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n202), .B2(new_n794), .C1(new_n1146), .C2(new_n890), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n386), .B(new_n1272), .C1(new_n814), .C2(new_n1142), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n812), .A2(G159), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n802), .A2(G137), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G128), .B2(new_n886), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n782), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n780), .B1(new_n203), .B2(new_n899), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n964), .A2(new_n837), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1278), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1263), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1193), .A2(new_n1199), .A3(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1288), .B2(new_n1011), .ZN(G381));
  NAND2_X1  g1089(.A1(new_n1261), .A2(new_n1203), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1290), .A2(G396), .A3(G393), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(G381), .A2(G384), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1072), .A2(new_n1074), .A3(G390), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(G407));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G343), .C2(new_n1290), .ZN(G409));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(G390), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1041), .B2(new_n1071), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1041), .A2(new_n1071), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(G390), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1302), .A2(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1297), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1010), .B(new_n1246), .C1(new_n1256), .C2(new_n1192), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1203), .A2(new_n1308), .A3(new_n1247), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n708), .A2(G213), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G378), .B2(new_n1259), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT60), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n736), .B(new_n1313), .C1(new_n1288), .C2(KEYINPUT60), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n901), .B(new_n875), .C1(new_n1314), .C2(new_n1285), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(new_n1288), .B2(KEYINPUT60), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n735), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(G384), .A3(new_n1286), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1307), .B1(new_n1312), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT57), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1246), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1192), .B1(new_n1183), .B2(new_n1200), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1322), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n735), .A3(new_n1257), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1203), .B1(new_n1326), .B2(new_n1247), .ZN(new_n1327));
  NOR4_X1   g1127(.A1(new_n1327), .A2(new_n1311), .A3(new_n1319), .A4(KEYINPUT62), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1321), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n708), .A2(G213), .A3(G2897), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1315), .A2(new_n1318), .A3(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1330), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1259), .A2(G378), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1311), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT61), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1306), .B1(new_n1329), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1333), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1340), .B(new_n1331), .C1(new_n1327), .C2(new_n1311), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1341), .A2(KEYINPUT63), .B1(new_n1312), .B2(new_n1320), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1305), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1320), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1296), .B1(new_n1339), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(KEYINPUT62), .B1(new_n1337), .B2(new_n1319), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1312), .A2(new_n1307), .A3(new_n1320), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1338), .A2(new_n1348), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1306), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1353), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1337), .A2(new_n1319), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1343), .B(new_n1344), .C1(new_n1354), .C2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1352), .A2(KEYINPUT126), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1347), .A2(new_n1357), .ZN(G405));
  NAND2_X1  g1158(.A1(new_n1320), .A2(KEYINPUT127), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1290), .A2(new_n1335), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1359), .B1(new_n1290), .B2(new_n1335), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1306), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1362), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1364), .A2(new_n1351), .A3(new_n1360), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1363), .A2(new_n1365), .ZN(G402));
endmodule


