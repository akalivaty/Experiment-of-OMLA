//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n640, new_n641, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n462), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n471), .B2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n475), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OR2_X1    g064(.A1(new_n462), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT68), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n462), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n493), .A2(new_n496), .B1(new_n484), .B2(G126), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n465), .A2(new_n500), .A3(G138), .A4(new_n462), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT70), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(KEYINPUT69), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n507), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G88), .B1(new_n518), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n512), .B2(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n521), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n515), .A2(G89), .ZN(new_n526));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n527), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT71), .B(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n515), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n521), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n507), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(G43), .A2(new_n521), .B1(new_n515), .B2(G81), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n507), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n546), .A2(new_n548), .A3(G651), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n510), .B1(KEYINPUT70), .B2(G651), .ZN(new_n559));
  INV_X1    g134(.A(G651), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT6), .B1(new_n560), .B2(KEYINPUT69), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n514), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  AND3_X1   g138(.A1(KEYINPUT73), .A2(G53), .A3(G543), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n558), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n564), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(KEYINPUT74), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n515), .A2(G91), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT75), .B1(new_n505), .B2(new_n506), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(new_n520), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(KEYINPUT5), .A2(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n574), .B1(new_n581), .B2(G65), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n573), .B1(new_n582), .B2(new_n560), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n572), .A2(new_n584), .ZN(G299));
  NAND2_X1  g160(.A1(G171), .A2(KEYINPUT76), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G301));
  NAND2_X1  g166(.A1(new_n521), .A2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n515), .A2(G87), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(new_n515), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n521), .A2(G48), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n507), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n607), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n599), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(G72), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n507), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(new_n614), .C1(new_n507), .C2(new_n615), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(G651), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n521), .A2(G47), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n515), .A2(G85), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(new_n521), .A2(G54), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n575), .B2(new_n580), .ZN(new_n629));
  AND2_X1   g204(.A1(G79), .A2(G543), .ZN(new_n630));
  OAI21_X1  g205(.A(G651), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(KEYINPUT10), .B1(new_n515), .B2(G92), .ZN(new_n632));
  AND4_X1   g207(.A1(KEYINPUT10), .A2(new_n562), .A3(G92), .A4(new_n527), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n627), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n590), .B2(G868), .ZN(G284));
  AOI21_X1  g211(.A(new_n635), .B1(new_n590), .B2(G868), .ZN(G321));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NOR2_X1   g213(.A1(G286), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n583), .B1(new_n567), .B2(new_n571), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n639), .B1(new_n641), .B2(new_n638), .ZN(G297));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n638), .ZN(G280));
  NOR2_X1   g218(.A1(new_n632), .A2(new_n633), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n631), .A2(new_n627), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(G860), .ZN(G148));
  NOR2_X1   g223(.A1(new_n634), .A2(G559), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  MUX2_X1   g225(.A(new_n551), .B(new_n650), .S(G868), .Z(G323));
  XNOR2_X1  g226(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g227(.A1(new_n484), .A2(G123), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n462), .A2(G111), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  INV_X1    g230(.A(G135), .ZN(new_n656));
  OAI221_X1 g231(.A(new_n653), .B1(new_n654), .B2(new_n655), .C1(new_n656), .C2(new_n466), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n465), .A2(new_n463), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT12), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT13), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n663), .ZN(G156));
  XNOR2_X1  g239(.A(G2427), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(KEYINPUT14), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2443), .B(G2446), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2451), .B(G2454), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1341), .B(G1348), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT85), .Z(new_n680));
  INV_X1    g255(.A(G14), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n678), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT86), .Z(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(G401));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  XOR2_X1   g261(.A(G2084), .B(G2090), .Z(new_n687));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(KEYINPUT17), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n688), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2100), .ZN(new_n693));
  XOR2_X1   g268(.A(G2072), .B(G2078), .Z(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n689), .B2(KEYINPUT18), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2096), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1971), .B(G1976), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n700), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(KEYINPUT87), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT20), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT88), .ZN(new_n711));
  XOR2_X1   g286(.A(G1981), .B(G1986), .Z(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n711), .B(new_n716), .ZN(G229));
  NAND2_X1  g292(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G1986), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G131), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G107), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G119), .B2(new_n484), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G25), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n722), .A2(G1986), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n723), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n719), .A2(G22), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G166), .B2(new_n719), .ZN(new_n739));
  INV_X1    g314(.A(G1971), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G23), .B(G288), .S(G16), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT33), .B(G1976), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT32), .B(G1981), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n719), .A2(G6), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n612), .B2(new_n719), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n741), .B(new_n744), .C1(new_n745), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n736), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n749), .A2(new_n737), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n718), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G32), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n484), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(new_n756), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G28), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT30), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(KEYINPUT30), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n766), .B(new_n772), .C1(new_n756), .C2(new_n658), .ZN(new_n773));
  NOR2_X1   g348(.A1(G171), .A2(new_n719), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G5), .B2(new_n719), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G1961), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n484), .A2(G128), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n462), .A2(G116), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  INV_X1    g355(.A(G140), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n778), .B1(new_n779), .B2(new_n780), .C1(new_n781), .C2(new_n466), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n756), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n756), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n756), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(G2078), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n773), .A2(new_n777), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(G286), .A2(G16), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n719), .A2(G21), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT24), .ZN(new_n800));
  INV_X1    g375(.A(G34), .ZN(new_n801));
  AOI21_X1  g376(.A(G29), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G160), .B2(new_n756), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n799), .A2(G1966), .B1(G2084), .B2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G1966), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n776), .A2(G1961), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(G2084), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT94), .Z(new_n809));
  NOR2_X1   g384(.A1(G4), .A2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT91), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n634), .B2(new_n719), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1348), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n795), .A2(new_n805), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n756), .A2(G33), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G139), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n466), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n465), .A2(G127), .ZN(new_n822));
  NAND2_X1  g397(.A1(G115), .A2(G2104), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n462), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n826), .B2(new_n756), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(G2072), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n719), .A2(G20), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT23), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n640), .B2(new_n719), .ZN(new_n831));
  INV_X1    g406(.A(G1956), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n719), .A2(G19), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT92), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n552), .B2(new_n719), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n756), .A2(G35), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT95), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G162), .B2(new_n756), .ZN(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n828), .A2(new_n833), .A3(new_n837), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n815), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT97), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n755), .A2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n755), .A2(new_n847), .ZN(G150));
  NAND2_X1  g424(.A1(new_n521), .A2(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n515), .A2(G93), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n507), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT98), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n551), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n547), .B(new_n548), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n543), .A4(new_n857), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT38), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n646), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n856), .A2(G860), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n870), .A2(new_n872), .ZN(G145));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n658), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n658), .B(KEYINPUT99), .ZN(new_n877));
  INV_X1    g452(.A(G160), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n488), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n876), .A2(new_n879), .A3(G162), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n731), .B(new_n661), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n480), .A2(G142), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n484), .A2(G130), .ZN(new_n890));
  OR2_X1    g465(.A1(G106), .A2(G2105), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n891), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n782), .B(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(G164), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(G164), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n763), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n905), .A2(new_n901), .A3(new_n762), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n904), .A2(new_n906), .A3(new_n825), .ZN(new_n907));
  INV_X1    g482(.A(new_n826), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n762), .B1(new_n905), .B2(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n763), .A3(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n887), .B(new_n898), .C1(new_n907), .C2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n897), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n887), .B1(new_n913), .B2(new_n895), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n896), .A2(KEYINPUT101), .A3(new_n897), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n826), .B1(new_n904), .B2(new_n906), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n909), .B(new_n910), .C1(new_n824), .C2(new_n821), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n886), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n881), .A2(new_n883), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(KEYINPUT102), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(KEYINPUT102), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g501(.A1(new_n721), .A2(G305), .ZN(new_n927));
  XNOR2_X1  g502(.A(G303), .B(G288), .ZN(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(new_n612), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n927), .B2(new_n929), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n931), .B2(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n650), .B(new_n864), .Z(new_n940));
  NAND3_X1  g515(.A1(G299), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n640), .B2(new_n634), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n941), .A2(new_n943), .B1(new_n640), .B2(new_n634), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n640), .B2(new_n634), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT104), .B1(G299), .B2(new_n646), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n640), .A2(new_n942), .A3(new_n634), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n941), .A2(new_n943), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n947), .ZN(new_n954));
  NAND2_X1  g529(.A1(G299), .A2(new_n646), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n572), .A2(new_n634), .A3(new_n584), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT41), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n945), .B1(new_n940), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n939), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n934), .A2(KEYINPUT106), .A3(new_n936), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n939), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g538(.A(G868), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(G868), .B2(new_n857), .ZN(G295));
  OAI21_X1  g540(.A(new_n964), .B1(G868), .B2(new_n857), .ZN(G331));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  NOR2_X1   g544(.A1(G168), .A2(G171), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n590), .B2(G168), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n864), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G286), .B1(new_n586), .B2(new_n589), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n863), .B(new_n861), .C1(new_n973), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n957), .B1(new_n950), .B2(KEYINPUT105), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n969), .B(new_n975), .C1(new_n976), .C2(new_n954), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n972), .A2(new_n974), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT107), .B1(new_n959), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n944), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n933), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n956), .A2(KEYINPUT41), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n943), .B2(new_n941), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n958), .B1(new_n984), .B2(new_n953), .ZN(new_n985));
  INV_X1    g560(.A(new_n954), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n969), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n959), .A2(KEYINPUT107), .A3(new_n978), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n932), .ZN(new_n991));
  INV_X1    g566(.A(new_n944), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n991), .A2(new_n930), .B1(new_n992), .B2(new_n975), .ZN(new_n993));
  AOI21_X1  g568(.A(G37), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n968), .B1(new_n982), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n993), .B1(new_n977), .B2(new_n979), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n947), .A2(new_n955), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT41), .B1(new_n952), .B2(new_n956), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(KEYINPUT108), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n944), .B2(KEYINPUT41), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n975), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n933), .B1(new_n1003), .B2(new_n981), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n997), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n967), .B1(new_n995), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n996), .A2(KEYINPUT109), .A3(new_n1004), .A4(new_n997), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1009), .A2(KEYINPUT43), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n982), .A2(new_n994), .A3(new_n968), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT44), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1007), .B1(new_n1011), .B2(new_n1013), .ZN(G397));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n503), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n471), .A2(new_n478), .ZN(new_n1019));
  INV_X1    g594(.A(new_n468), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(G40), .A3(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(G1996), .A3(new_n762), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1024));
  XNOR2_X1  g599(.A(new_n782), .B(new_n787), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(G1996), .B2(new_n762), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1022), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n731), .B(new_n733), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OR3_X1    g605(.A1(G290), .A2(new_n1028), .A3(G1986), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G290), .A2(G1986), .A3(new_n1022), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT110), .Z(new_n1034));
  NOR2_X1   g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  INV_X1    g611(.A(G40), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n1037), .B(new_n468), .C1(new_n471), .C2(new_n478), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1018), .A2(new_n1038), .A3(new_n789), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1038), .A3(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT125), .B(G1961), .Z(new_n1046));
  AOI22_X1  g621(.A1(new_n1036), .A2(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1018), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G301), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1045), .B2(G2084), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n1021), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1056), .A2(KEYINPUT118), .A3(new_n1057), .A4(new_n1044), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1048), .A2(new_n806), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(G286), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1054), .A2(new_n1058), .A3(G168), .A4(new_n1059), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G8), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1062), .A2(new_n1065), .A3(G8), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1052), .B1(new_n1068), .B2(KEYINPUT62), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1045), .A2(KEYINPUT115), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1042), .A2(new_n1038), .A3(new_n1072), .A4(new_n1044), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n841), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1048), .A2(new_n740), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1070), .B1(new_n1076), .B2(KEYINPUT116), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1078), .A3(new_n1075), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G303), .A2(G8), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1081), .B(KEYINPUT55), .Z(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1021), .B2(new_n1016), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  OR2_X1    g662(.A1(G288), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT52), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n1091));
  AOI211_X1 g666(.A(G1981), .B(new_n599), .C1(new_n608), .C2(new_n611), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n606), .A2(new_n607), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n598), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n612), .A2(new_n1093), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1095), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(KEYINPUT49), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1099), .A3(new_n1086), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1056), .A2(new_n841), .A3(new_n1044), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1070), .B1(new_n1101), .B2(new_n1075), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1082), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1086), .A2(new_n1088), .A3(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1090), .A2(new_n1100), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1082), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1060), .A2(G286), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(new_n1062), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1066), .B1(new_n1111), .B2(KEYINPUT51), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1069), .A2(new_n1083), .A3(new_n1109), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1045), .A2(new_n832), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1018), .A2(new_n1038), .A3(new_n1040), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n569), .B2(new_n570), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n584), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n640), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1121), .B(new_n1125), .C1(new_n640), .C2(new_n1122), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT121), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1124), .A2(new_n1130), .A3(new_n1126), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1119), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1348), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1021), .A2(new_n1016), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1045), .A2(new_n1133), .B1(new_n1134), .B2(new_n787), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n634), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1127), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1138));
  AND4_X1   g713(.A1(new_n1124), .A2(new_n1118), .A3(new_n1126), .A4(new_n1116), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1124), .A2(new_n1126), .B1(new_n1118), .B2(new_n1116), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n646), .B2(KEYINPUT124), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n646), .A2(KEYINPUT124), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1135), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1135), .B2(new_n1143), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT58), .B(G1341), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1048), .A2(G1996), .B1(new_n1134), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n552), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1141), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1127), .A2(KEYINPUT61), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1132), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1137), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1041), .A2(new_n1036), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n477), .A2(G2105), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n468), .A2(new_n1037), .A3(new_n1049), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1018), .A2(new_n1159), .A3(new_n1040), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G171), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1047), .A2(G301), .A3(new_n1050), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(KEYINPUT54), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1163), .A2(new_n590), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1167), .A2(new_n1051), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1168), .B2(KEYINPUT54), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1112), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1157), .A2(new_n1170), .A3(new_n1083), .A4(new_n1109), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1090), .A2(new_n1105), .A3(new_n1100), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1103), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G288), .A2(G1976), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT114), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1100), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1097), .B(KEYINPUT113), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1172), .A2(new_n1173), .B1(new_n1178), .B2(new_n1086), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1115), .A2(new_n1171), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT63), .B1(new_n1102), .B2(new_n1082), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1060), .A2(G8), .A3(G168), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1172), .A2(new_n1181), .A3(new_n1103), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1184), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT119), .B1(new_n1186), .B2(new_n1106), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1183), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1083), .A2(new_n1109), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1188), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1035), .B1(new_n1180), .B2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1027), .A2(new_n733), .A3(new_n726), .A4(new_n730), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n782), .A2(G2067), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1028), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1028), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT46), .B1(new_n1028), .B2(G1996), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1025), .A2(new_n763), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1197), .A2(new_n1198), .B1(new_n1022), .B2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT47), .Z(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT127), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1031), .B(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1030), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1196), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1193), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g782(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1209));
  AOI21_X1  g783(.A(new_n1209), .B1(new_n682), .B2(new_n684), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n1210), .B(new_n925), .C1(new_n995), .C2(new_n1006), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


