//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT66), .B(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n463), .C1(new_n469), .C2(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n468), .B1(new_n472), .B2(new_n461), .ZN(G160));
  OAI211_X1 g048(.A(new_n461), .B(new_n463), .C1(new_n469), .C2(new_n462), .ZN(new_n474));
  INV_X1    g049(.A(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G2105), .A3(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n478), .B1(G124), .B2(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT4), .B1(new_n474), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n482), .A2(G138), .A3(new_n461), .A4(new_n463), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .A3(KEYINPUT4), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n463), .A2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(new_n461), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n484), .A2(G126), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT69), .B1(new_n505), .B2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G62), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(new_n520), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NOR2_X1   g100(.A1(new_n512), .A2(new_n515), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n512), .A2(new_n519), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(G90), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n526), .A2(G43), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT71), .B(G81), .Z(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n519), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n544), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  XOR2_X1   g129(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n526), .A2(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n526), .A2(KEYINPUT9), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n519), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n528), .A2(G91), .B1(new_n565), .B2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n526), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n528), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n520), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n508), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n526), .A2(G48), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n526), .A2(KEYINPUT73), .A3(G48), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n522), .ZN(G305));
  AOI22_X1  g157(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  AOI22_X1  g160(.A1(G47), .A2(new_n526), .B1(new_n528), .B2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n528), .A2(new_n588), .A3(G92), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n528), .B2(G92), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n519), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n526), .A2(G54), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G171), .B2(new_n597), .ZN(G284));
  OAI21_X1  g174(.A(new_n598), .B1(G171), .B2(new_n597), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(new_n596), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g186(.A1(new_n492), .A2(new_n469), .A3(new_n461), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n461), .A2(G111), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT75), .Z(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n484), .A2(G123), .ZN(new_n619));
  INV_X1    g194(.A(new_n474), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G135), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2435), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2438), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2451), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT77), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n643), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n640), .B(KEYINPUT78), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n640), .B(KEYINPUT17), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(new_n647), .ZN(new_n650));
  OAI221_X1 g225(.A(new_n646), .B1(new_n647), .B2(new_n648), .C1(new_n650), .C2(new_n644), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2100), .Z(G227));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  AOI22_X1  g237(.A1(new_n660), .A2(new_n661), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n657), .A2(new_n662), .A3(new_n659), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n663), .B(new_n664), .C1(new_n661), .C2(new_n660), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(G1986), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT22), .B(G1981), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  NAND2_X1  g247(.A1(new_n484), .A2(G119), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n620), .A2(G131), .ZN(new_n674));
  NOR2_X1   g249(.A1(G95), .A2(G2105), .ZN(new_n675));
  OAI21_X1  g250(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  MUX2_X1   g254(.A(G25), .B(new_n679), .S(G29), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT35), .B(G1991), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT82), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n683), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G1971), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n694), .B1(new_n693), .B2(new_n697), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n682), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G24), .ZN(new_n701));
  XOR2_X1   g276(.A(G290), .B(KEYINPUT81), .Z(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n700), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(G29), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT25), .Z(new_n713));
  INV_X1    g288(.A(G139), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n713), .B1(new_n474), .B2(new_n714), .C1(new_n715), .C2(new_n461), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G164), .A2(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G27), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G34), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G160), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n731), .A2(new_n732), .B1(new_n718), .B2(new_n719), .ZN(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G32), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n484), .A2(G129), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n482), .A2(G141), .A3(new_n463), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n469), .A2(G105), .ZN(new_n737));
  AOI21_X1  g312(.A(G2105), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT85), .B(KEYINPUT26), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n735), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  OAI211_X1 g319(.A(new_n724), .B(new_n733), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n683), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n551), .B2(new_n683), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1341), .Z(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n722), .B2(new_n723), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n717), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n622), .B2(new_n717), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT87), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n745), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n732), .B2(new_n731), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n717), .A2(G26), .ZN(new_n758));
  INV_X1    g333(.A(G140), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n484), .A2(G128), .ZN(new_n761));
  NOR2_X1   g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT83), .B1(new_n474), .B2(new_n759), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n760), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(new_n717), .ZN(new_n769));
  MUX2_X1   g344(.A(new_n758), .B(new_n769), .S(KEYINPUT28), .Z(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2067), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n683), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n605), .B2(new_n683), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n683), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n683), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT86), .B(G1966), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT88), .B(KEYINPUT23), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n683), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n602), .B2(new_n683), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n743), .B2(new_n744), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n771), .A2(new_n775), .A3(new_n779), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n757), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n710), .A2(new_n720), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n717), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n717), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT29), .Z(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n683), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n683), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n788), .A2(new_n793), .A3(new_n798), .ZN(G311));
  AND2_X1   g374(.A1(new_n710), .A2(new_n787), .ZN(new_n800));
  INV_X1    g375(.A(new_n793), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n800), .A2(new_n801), .A3(new_n797), .A4(new_n720), .ZN(G150));
  NAND2_X1  g377(.A1(new_n528), .A2(G93), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT89), .B(G55), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n526), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(G80), .A2(G543), .ZN(new_n806));
  INV_X1    g381(.A(G67), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n519), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G651), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n803), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n803), .A2(new_n805), .A3(KEYINPUT91), .A4(new_n809), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G860), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NOR2_X1   g391(.A1(new_n596), .A2(new_n606), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n551), .B1(new_n812), .B2(new_n813), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n551), .A2(new_n810), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT90), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(KEYINPUT90), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n816), .B1(new_n825), .B2(G860), .ZN(G145));
  INV_X1    g401(.A(KEYINPUT93), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n716), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n679), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n484), .A2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n620), .A2(G142), .ZN(new_n831));
  NOR2_X1   g406(.A1(G106), .A2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n829), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n622), .B(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G162), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n613), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n835), .B(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n490), .A2(KEYINPUT68), .A3(KEYINPUT4), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT68), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n840), .A2(new_n841), .A3(new_n494), .ZN(new_n842));
  INV_X1    g417(.A(new_n502), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT92), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n496), .A2(new_n845), .A3(new_n502), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n767), .ZN(new_n848));
  INV_X1    g423(.A(new_n742), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n827), .B2(new_n716), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n839), .A2(new_n851), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g431(.A(G166), .B(new_n685), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(G305), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(G305), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G290), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(G290), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT42), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n596), .B(G299), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT94), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n596), .A2(new_n602), .A3(KEYINPUT94), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(KEYINPUT41), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n868), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT95), .Z(new_n874));
  AND2_X1   g449(.A1(new_n822), .A2(new_n823), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n608), .ZN(new_n876));
  MUX2_X1   g451(.A(new_n872), .B(new_n874), .S(new_n876), .Z(new_n877));
  AOI21_X1  g452(.A(new_n865), .B1(new_n877), .B2(KEYINPUT96), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(KEYINPUT96), .B2(new_n877), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n877), .A2(KEYINPUT96), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n597), .B1(new_n880), .B2(new_n865), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT97), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n879), .A2(new_n881), .B1(new_n597), .B2(new_n814), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n884), .B2(KEYINPUT97), .ZN(G295));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(KEYINPUT97), .ZN(G331));
  AND3_X1   g461(.A1(new_n862), .A2(KEYINPUT100), .A3(new_n863), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT100), .B1(new_n862), .B2(new_n863), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n866), .A2(new_n870), .ZN(new_n890));
  XNOR2_X1  g465(.A(G301), .B(G286), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n824), .B(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n890), .B(new_n892), .C1(new_n870), .C2(new_n873), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT99), .B1(new_n875), .B2(new_n891), .ZN(new_n894));
  INV_X1    g469(.A(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT98), .B1(new_n895), .B2(new_n824), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n875), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n895), .A2(new_n824), .A3(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n894), .A2(new_n896), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n874), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n889), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n872), .ZN(new_n904));
  INV_X1    g479(.A(new_n873), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n901), .A2(new_n904), .B1(new_n892), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(G37), .B1(new_n906), .B2(new_n864), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(KEYINPUT43), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n889), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT43), .B1(new_n910), .B2(new_n907), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT44), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n906), .A2(new_n864), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n853), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n887), .A2(new_n888), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n906), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT101), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n903), .A2(new_n919), .A3(new_n907), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(KEYINPUT43), .C1(new_n914), .C2(new_n916), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n912), .B1(new_n924), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n496), .A2(new_n845), .A3(new_n502), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n845), .B1(new_n496), .B2(new_n502), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  XOR2_X1   g505(.A(KEYINPUT102), .B(G40), .Z(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(G160), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  AOI21_X1  g509(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n935));
  NOR4_X1   g510(.A1(new_n935), .A2(KEYINPUT103), .A3(new_n468), .A4(new_n931), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n930), .A3(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT104), .Z(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(G1986), .A3(G290), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n704), .A3(new_n861), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT105), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n767), .B(G2067), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT106), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT107), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n940), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n742), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n679), .B(new_n681), .Z(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT108), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n940), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n948), .A2(new_n950), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n944), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(G1384), .C1(new_n496), .C2(new_n502), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n792), .B(new_n938), .C1(new_n960), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT45), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(G160), .B2(new_n932), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n936), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n926), .B1(new_n842), .B2(new_n843), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n930), .ZN(new_n970));
  AOI21_X1  g545(.A(G1971), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G303), .A2(G8), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT55), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT109), .B(G86), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n580), .B1(new_n522), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G1981), .ZN(new_n981));
  INV_X1    g556(.A(G1981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n580), .B(new_n982), .C1(new_n581), .C2(new_n522), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(KEYINPUT49), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n983), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n969), .A2(new_n968), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n973), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n981), .A2(new_n991), .A3(new_n983), .A4(KEYINPUT49), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n985), .A2(new_n988), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n990), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT52), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n995), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n990), .B(new_n998), .C1(new_n995), .C2(G288), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n983), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G288), .A2(G1976), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT111), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1001), .B1(new_n993), .B2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n978), .A2(new_n1000), .B1(new_n1004), .B2(new_n994), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n964), .B2(new_n971), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n938), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n844), .B2(new_n846), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1010));
  OAI211_X1 g585(.A(KEYINPUT112), .B(new_n963), .C1(new_n1010), .C2(G1971), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1011), .A3(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n976), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1000), .B1(new_n977), .B2(new_n974), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n969), .A2(new_n930), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n778), .B1(new_n1016), .B2(new_n1008), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n732), .B(new_n938), .C1(new_n960), .C2(new_n962), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(G168), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT51), .ZN(new_n1021));
  AOI21_X1  g596(.A(G168), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1019), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1012), .A2(new_n1027), .A3(new_n976), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1014), .A2(new_n1015), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n965), .A2(new_n970), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(G2078), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1016), .A2(new_n1008), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT53), .A3(new_n723), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n938), .B1(new_n960), .B2(new_n962), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n796), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1038), .A2(KEYINPUT120), .A3(G171), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT120), .B1(new_n1038), .B2(G171), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1030), .A2(KEYINPUT123), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1029), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1030), .A2(KEYINPUT123), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1005), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n929), .A2(new_n930), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G160), .A2(G40), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT53), .B(new_n723), .C1(new_n1046), .C2(KEYINPUT121), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(KEYINPUT121), .B2(new_n1046), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n965), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1033), .A2(new_n1037), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G171), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1033), .A2(new_n1035), .A3(G301), .A4(new_n1037), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(KEYINPUT54), .A3(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1014), .A2(new_n1015), .A3(new_n1028), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1036), .A2(new_n774), .ZN(new_n1057));
  INV_X1    g632(.A(new_n989), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(G2067), .B2(new_n1058), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1059), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT61), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1036), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n565), .A2(G651), .ZN(new_n1065));
  INV_X1    g640(.A(G91), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n522), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n566), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(new_n561), .A4(new_n562), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n1071), .B2(KEYINPUT115), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n602), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(KEYINPUT57), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n965), .A2(new_n970), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1064), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1064), .B2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1062), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1064), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(KEYINPUT119), .B2(new_n1061), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1060), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT58), .B(G1341), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1032), .A2(G1996), .B1(new_n989), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(KEYINPUT118), .A3(new_n551), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT117), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1088), .A3(new_n551), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(KEYINPUT59), .A3(new_n1089), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1059), .A2(new_n605), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1059), .A2(new_n605), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1086), .A2(KEYINPUT117), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1083), .A2(new_n1090), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1079), .B1(new_n1091), .B2(new_n1081), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1050), .A2(G171), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1039), .A2(new_n1040), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1101), .B2(KEYINPUT54), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1040), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1038), .A2(KEYINPUT120), .A3(G171), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT122), .B(new_n1103), .C1(new_n1106), .C2(new_n1100), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1056), .A2(new_n1098), .A3(new_n1102), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1044), .A2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n973), .B(G286), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1014), .A2(new_n1015), .A3(new_n1028), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n976), .B1(new_n972), .B2(new_n973), .ZN(new_n1116));
  AND4_X1   g691(.A1(KEYINPUT63), .A2(new_n1015), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n958), .B1(new_n1109), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT48), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT48), .A3(new_n1121), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1126), .A3(new_n957), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n679), .A2(new_n681), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n948), .A2(new_n950), .A3(new_n953), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(G2067), .B2(new_n767), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n940), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n940), .A2(new_n951), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT46), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n946), .A2(new_n849), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n940), .A2(new_n1137), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n940), .A2(KEYINPUT124), .A3(KEYINPUT46), .A4(new_n951), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT47), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT47), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1145), .A3(new_n1142), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1132), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1119), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g723(.A1(G401), .A2(G227), .ZN(new_n1150));
  AND2_X1   g724(.A1(new_n855), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n923), .A2(new_n1151), .A3(new_n459), .A4(new_n671), .ZN(G225));
  INV_X1    g726(.A(G225), .ZN(G308));
endmodule


