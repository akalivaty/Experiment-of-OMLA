//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1112,
    new_n1113, new_n1114;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n460), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n460), .B2(G112), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND4_X1  g056(.A1(new_n470), .A2(new_n472), .A3(G126), .A4(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n461), .A2(new_n484), .A3(G126), .A4(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n460), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n461), .A2(new_n489), .A3(G138), .A4(new_n460), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(new_n460), .B2(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n486), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(G75), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n506), .B(KEYINPUT69), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n500), .A2(new_n502), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G166));
  NOR2_X1   g094(.A1(new_n509), .A2(new_n510), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n499), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n511), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n522), .B(new_n524), .C1(new_n525), .C2(new_n503), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G168));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n512), .A2(new_n530), .B1(new_n514), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n532), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n512), .A2(new_n538), .B1(new_n514), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n534), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n545), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n511), .A2(KEYINPUT71), .A3(G543), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n521), .A2(KEYINPUT71), .A3(KEYINPUT9), .A4(G53), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT72), .ZN(new_n556));
  INV_X1    g131(.A(new_n512), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n503), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n557), .A2(G91), .B1(G651), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n553), .A2(new_n562), .A3(new_n554), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n556), .A2(new_n561), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  XNOR2_X1  g140(.A(new_n518), .B(KEYINPUT73), .ZN(G303));
  NAND2_X1  g141(.A1(new_n521), .A2(G49), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT74), .Z(new_n568));
  OR2_X1    g143(.A1(new_n508), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(G87), .A2(new_n557), .B1(new_n569), .B2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n512), .A2(new_n572), .B1(new_n514), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n534), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n534), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n557), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n521), .A2(G47), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(KEYINPUT75), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(G290));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n503), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT10), .B1(new_n512), .B2(new_n586), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G171), .B2(new_n594), .ZN(G284));
  OAI21_X1  g171(.A(new_n595), .B1(G171), .B2(new_n594), .ZN(G321));
  NAND2_X1  g172(.A1(G299), .A2(new_n594), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n594), .B2(G168), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(new_n594), .B2(G168), .ZN(G280));
  INV_X1    g175(.A(new_n593), .ZN(new_n601));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G860), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT76), .ZN(G148));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(KEYINPUT77), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n543), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n474), .A2(G123), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n476), .A2(G135), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT79), .ZN(new_n614));
  NOR2_X1   g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n612), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n476), .A2(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2435), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2438), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  NOR3_X1   g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(KEYINPUT83), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(KEYINPUT17), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n644), .C1(new_n642), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n642), .A2(new_n651), .A3(new_n643), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT86), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  INV_X1    g244(.A(new_n660), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n662), .A2(new_n663), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n670), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n669), .B(new_n673), .C1(new_n670), .C2(new_n672), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n568), .A2(new_n570), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT33), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n682), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n682), .A2(G6), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n577), .B2(new_n682), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n688), .A2(new_n692), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n698));
  OR2_X1    g273(.A1(G16), .A2(G24), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G290), .B2(new_n682), .ZN(new_n700));
  INV_X1    g275(.A(G1986), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(KEYINPUT91), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n474), .A2(G119), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n476), .A2(G131), .ZN(new_n709));
  OR2_X1    g284(.A1(G95), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(new_n706), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n707), .B(new_n714), .S(KEYINPUT88), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT89), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n705), .B(new_n718), .C1(new_n701), .C2(new_n700), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n682), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n682), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G1966), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT92), .B1(G4), .B2(G16), .ZN(new_n725));
  OR3_X1    g300(.A1(KEYINPUT92), .A2(G4), .A3(G16), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(new_n593), .C2(new_n682), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1348), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n476), .A2(G140), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n461), .A2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G128), .ZN(new_n733));
  NOR2_X1   g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n706), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n739), .A2(G2067), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(G2067), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n724), .B(new_n728), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT100), .B1(G5), .B2(G16), .ZN(new_n745));
  OR3_X1    g320(.A1(KEYINPUT100), .A2(G5), .A3(G16), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n745), .B(new_n746), .C1(G301), .C2(new_n682), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1961), .Z(new_n748));
  NAND2_X1  g323(.A1(G164), .A2(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(G27), .A2(G29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(G2078), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n682), .A2(KEYINPUT23), .A3(G20), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n755));
  INV_X1    g330(.A(G20), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G299), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n754), .B(new_n757), .C1(new_n758), .C2(new_n682), .ZN(new_n759));
  INV_X1    g334(.A(G1956), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n706), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n706), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT29), .Z(new_n765));
  OAI211_X1 g340(.A(new_n753), .B(new_n761), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n618), .A2(G29), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n744), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G16), .A2(G19), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n543), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT93), .B(G1341), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(KEYINPUT24), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(KEYINPUT24), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n706), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G160), .B2(new_n706), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(G2084), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n765), .A2(new_n762), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT25), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n476), .A2(G139), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n783), .C1(new_n460), .C2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G2072), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G11), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT30), .B(G28), .Z(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n777), .B2(G2084), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n768), .A2(new_n779), .A3(new_n780), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G32), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT98), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT26), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT97), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n476), .A2(G141), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n474), .A2(G129), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n795), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT27), .B(G1996), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n723), .A2(G1966), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT99), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n794), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G2078), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n751), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n812), .A2(KEYINPUT101), .A3(new_n814), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n721), .B1(new_n817), .B2(new_n818), .ZN(G311));
  INV_X1    g394(.A(new_n721), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n812), .A2(KEYINPUT101), .A3(new_n814), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT101), .B1(new_n812), .B2(new_n814), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(G150));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n512), .A2(new_n824), .B1(new_n514), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n534), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT103), .B(G860), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  INV_X1    g408(.A(new_n829), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n543), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n829), .B1(new_n542), .B2(new_n540), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n593), .A2(new_n602), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT102), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n833), .B1(new_n843), .B2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(new_n805), .B(new_n496), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(new_n737), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n737), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n785), .B(KEYINPUT104), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G130), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n732), .A2(KEYINPUT105), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT105), .B1(new_n732), .B2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n476), .A2(G142), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n713), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT106), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n621), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n785), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n847), .B2(new_n848), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n851), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT107), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n618), .B(G160), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n851), .A2(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(new_n861), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n865), .A3(KEYINPUT107), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n865), .A3(new_n868), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g452(.A1(new_n834), .A2(new_n594), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n837), .B(new_n605), .ZN(new_n879));
  XNOR2_X1  g454(.A(G299), .B(new_n593), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(KEYINPUT41), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n879), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(G288), .B(new_n577), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n518), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G290), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n884), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n878), .B1(new_n888), .B2(new_n594), .ZN(G295));
  OAI21_X1  g464(.A(new_n878), .B1(new_n888), .B2(new_n594), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n891));
  OAI21_X1  g466(.A(G286), .B1(new_n891), .B2(G171), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n835), .A3(new_n836), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n837), .B(G286), .C1(new_n891), .C2(G171), .ZN(new_n894));
  NOR2_X1   g469(.A1(G301), .A2(KEYINPUT109), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n893), .B2(new_n894), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n896), .A2(new_n882), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n880), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(new_n887), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n901), .A3(G37), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n905), .B(KEYINPUT44), .C1(new_n906), .C2(new_n902), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n902), .A2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n904), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n910), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g486(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n912));
  INV_X1    g487(.A(G1384), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n496), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G160), .A2(G40), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n737), .B(G2067), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n805), .A2(G1996), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n805), .A2(G1996), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n712), .B(new_n717), .Z(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(G290), .A2(G1986), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n917), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT48), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n917), .B1(new_n918), .B2(new_n805), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n915), .A2(G1996), .A3(new_n916), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(KEYINPUT46), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(KEYINPUT46), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT126), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT47), .Z(new_n934));
  NAND2_X1  g509(.A1(new_n713), .A2(new_n717), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n921), .A2(new_n935), .B1(G2067), .B2(new_n737), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n927), .B(new_n934), .C1(new_n917), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n496), .A2(new_n913), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n939));
  INV_X1    g514(.A(new_n912), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n494), .B1(new_n483), .B2(new_n485), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n491), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT112), .B1(new_n943), .B2(new_n912), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n464), .A2(new_n467), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(KEYINPUT45), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n941), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n938), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(KEYINPUT50), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n916), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n948), .A2(new_n691), .B1(new_n952), .B2(new_n762), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n956));
  NAND3_X1  g531(.A1(G303), .A2(new_n956), .A3(G8), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT73), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n507), .B2(new_n517), .ZN(new_n960));
  OAI21_X1  g535(.A(G8), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT55), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n955), .A2(new_n963), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1981), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n577), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n968), .B2(new_n577), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n943), .A2(new_n946), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n971), .B(KEYINPUT49), .C1(new_n968), .C2(new_n577), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n684), .B2(G1976), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n980), .B(new_n981), .C1(G1976), .C2(new_n684), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2084), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n943), .A2(KEYINPUT50), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n949), .B(G1384), .C1(new_n942), .C2(new_n491), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n946), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n916), .B1(new_n943), .B2(new_n912), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n943), .A2(KEYINPUT45), .ZN(new_n991));
  AOI21_X1  g566(.A(G1966), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(G8), .B(G168), .C1(new_n989), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n967), .A2(new_n984), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n964), .B1(new_n966), .B2(KEYINPUT114), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n955), .A2(new_n997), .A3(new_n963), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n984), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n993), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n995), .B1(new_n1000), .B2(KEYINPUT63), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n979), .A2(new_n1002), .A3(new_n684), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n976), .B1(new_n1003), .B2(new_n971), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n984), .B2(new_n966), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT120), .B1(new_n989), .B2(new_n992), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n946), .B1(new_n938), .B2(new_n940), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n943), .A2(KEYINPUT45), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1008), .B(new_n988), .C1(new_n1011), .C2(G1966), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G168), .A2(new_n954), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1007), .A2(KEYINPUT121), .A3(G8), .A4(new_n1012), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT51), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n993), .A2(new_n1021), .A3(new_n1017), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(KEYINPUT122), .A3(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1007), .A2(new_n1016), .A3(new_n1012), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1016), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(new_n1018), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n948), .B2(G2078), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n952), .A2(G1961), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1011), .A2(KEYINPUT53), .A3(new_n813), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G171), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1023), .A2(new_n1028), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI22_X1  g618(.A1(new_n948), .A2(new_n1043), .B1(new_n952), .B2(G1956), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n555), .A2(KEYINPUT57), .ZN(new_n1045));
  AOI22_X1  g620(.A1(G299), .A2(KEYINPUT57), .B1(new_n561), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n952), .A2(G1348), .B1(G2067), .B2(new_n975), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT116), .A3(new_n601), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n975), .A2(G2067), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n946), .B1(new_n986), .B2(new_n987), .ZN(new_n1053));
  INV_X1    g628(.A(G1348), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1051), .B1(new_n1055), .B2(new_n593), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1048), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n916), .B1(new_n914), .B2(new_n939), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(new_n947), .A3(new_n944), .A4(new_n1042), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1053), .A2(new_n760), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1046), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT115), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1060), .A3(new_n1046), .A4(new_n1063), .ZN(new_n1064));
  AND4_X1   g639(.A1(new_n1041), .A2(new_n1057), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1041), .B1(new_n1066), .B2(new_n1057), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1044), .A2(KEYINPUT118), .A3(new_n1047), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1062), .A3(new_n1064), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT61), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1055), .A2(KEYINPUT60), .B1(new_n1075), .B2(new_n601), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1049), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n593), .B(new_n1075), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1078), .A2(new_n1080), .B1(new_n1061), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n975), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n948), .B2(G1996), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n543), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT59), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1074), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1029), .B(G2078), .C1(new_n916), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n915), .A3(new_n947), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1030), .A2(new_n1031), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1036), .B(new_n1037), .C1(G171), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1033), .A2(G171), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1094), .B2(G171), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1095), .A2(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1089), .A2(new_n1099), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1038), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1040), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n999), .B(KEYINPUT125), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1006), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(G290), .A2(G1986), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n917), .B1(new_n1106), .B2(new_n924), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n923), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1108), .B(KEYINPUT111), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n937), .B1(new_n1105), .B2(new_n1109), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g685(.A(G229), .B1(new_n874), .B2(new_n875), .ZN(new_n1112));
  NAND3_X1  g686(.A1(new_n638), .A2(G319), .A3(new_n656), .ZN(new_n1113));
  XNOR2_X1  g687(.A(new_n1113), .B(KEYINPUT127), .ZN(new_n1114));
  OAI211_X1 g688(.A(new_n1112), .B(new_n1114), .C1(new_n908), .C2(new_n909), .ZN(G225));
  INV_X1    g689(.A(G225), .ZN(G308));
endmodule


