//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT64), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT66), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n466), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n468), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n476), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n463), .B1(new_n469), .B2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n466), .A2(new_n472), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n492), .B2(KEYINPUT68), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n476), .B2(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n463), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n483), .A2(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT69), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(new_n518), .A3(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G88), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n520), .A2(new_n524), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G51), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n513), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n521), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  INV_X1    g117(.A(G77), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n527), .A2(new_n542), .B1(new_n543), .B2(new_n514), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI221_X1 g121(.A(KEYINPUT70), .B1(new_n543), .B2(new_n514), .C1(new_n527), .C2(new_n542), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G651), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT71), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT72), .B(G90), .Z(new_n550));
  AOI22_X1  g125(.A1(new_n528), .A2(new_n550), .B1(new_n515), .B2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n523), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n528), .A2(G81), .ZN(new_n556));
  AOI211_X1 g131(.A(new_n555), .B(new_n556), .C1(G43), .C2(new_n515), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  AND2_X1   g138(.A1(new_n521), .A2(G65), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT74), .Z(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n528), .A2(G91), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n515), .A2(G53), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT73), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n515), .A2(new_n572), .A3(G53), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n569), .B(new_n574), .C1(KEYINPUT9), .C2(new_n571), .ZN(G299));
  OAI21_X1  g150(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT75), .Z(new_n577));
  AOI22_X1  g152(.A1(G87), .A2(new_n528), .B1(new_n515), .B2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  AOI22_X1  g154(.A1(G86), .A2(new_n528), .B1(new_n515), .B2(G48), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n584), .B(G61), .C1(new_n525), .C2(new_n526), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n584), .B1(new_n521), .B2(G61), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n581), .B(G651), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT76), .B1(new_n527), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(new_n585), .A3(new_n583), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n581), .B1(new_n592), .B2(G651), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n580), .B1(new_n589), .B2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(G85), .A2(new_n528), .B1(new_n515), .B2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n523), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n528), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n527), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n515), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n605), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n605), .B2(G168), .ZN(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT79), .B(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(G860), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g190(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n466), .A2(new_n472), .ZN(new_n620));
  NOR3_X1   g195(.A1(new_n620), .A2(new_n468), .A3(G2105), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT82), .B(G2100), .Z(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n476), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n463), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n642), .B2(new_n643), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n639), .B(new_n645), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n647), .ZN(G401));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(G2072), .A2(G2078), .ZN(new_n662));
  OAI22_X1  g237(.A1(new_n656), .A2(new_n660), .B1(new_n444), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  INV_X1    g250(.A(new_n669), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n673), .C2(new_n677), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  OAI21_X1  g260(.A(KEYINPUT93), .B1(G29), .B2(G32), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n476), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n483), .A2(G129), .ZN(new_n688));
  NAND3_X1  g263(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT26), .Z(new_n690));
  AND3_X1   g265(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G29), .ZN(new_n692));
  MUX2_X1   g267(.A(KEYINPUT93), .B(new_n686), .S(new_n692), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT27), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT94), .B(G28), .Z(new_n696));
  AOI21_X1  g271(.A(G29), .B1(new_n696), .B2(KEYINPUT30), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(KEYINPUT30), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G11), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n698), .B(new_n699), .C1(new_n633), .C2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NOR2_X1   g277(.A1(G168), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n702), .B2(G21), .ZN(new_n704));
  INV_X1    g279(.A(G1966), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n695), .B(new_n706), .C1(new_n705), .C2(new_n704), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n612), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G4), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1348), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT86), .B(G16), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G19), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n557), .B2(new_n713), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(G1341), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G35), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n700), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT29), .B(G2090), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n709), .A2(new_n710), .ZN(new_n723));
  NOR4_X1   g298(.A1(new_n707), .A2(new_n717), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G299), .A2(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n712), .A2(G20), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT97), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1956), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n700), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n700), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2078), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n700), .B1(new_n735), .B2(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G34), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G160), .B2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2084), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n700), .A2(G33), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT25), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n466), .A2(new_n472), .A3(G127), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n463), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n742), .B(new_n745), .C1(G139), .C2(new_n476), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n740), .B1(new_n746), .B2(new_n700), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(new_n442), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n724), .A2(new_n734), .A3(new_n739), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n700), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n483), .A2(G128), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT91), .Z(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G116), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G2105), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G140), .B2(new_n476), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n758), .A2(KEYINPUT92), .A3(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(KEYINPUT92), .B1(new_n758), .B2(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n751), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n702), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n702), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n738), .A2(G2084), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  NAND4_X1  g344(.A1(new_n763), .A2(new_n766), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n749), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n702), .A2(G23), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G288), .B2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n713), .A2(G22), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n713), .ZN(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G6), .B(G305), .S(G16), .Z(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT32), .B(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT34), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n774), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(KEYINPUT88), .B(KEYINPUT34), .C1(new_n784), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n483), .A2(G119), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n476), .A2(G131), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n463), .A2(G107), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G25), .B(new_n797), .S(G29), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n712), .A2(G24), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT87), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G290), .B2(new_n713), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1986), .Z(new_n805));
  AOI211_X1 g380(.A(new_n801), .B(new_n805), .C1(new_n788), .C2(new_n789), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n773), .B1(new_n792), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n792), .A2(new_n806), .A3(new_n773), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n808), .A2(KEYINPUT89), .A3(KEYINPUT36), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n811));
  INV_X1    g386(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n807), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n772), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(G311));
  INV_X1    g391(.A(new_n814), .ZN(G150));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n527), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n523), .B1(new_n820), .B2(KEYINPUT99), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(KEYINPUT99), .B2(new_n820), .ZN(new_n822));
  AOI22_X1  g397(.A1(G93), .A2(new_n528), .B1(new_n515), .B2(G55), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n612), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n557), .B(new_n824), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT100), .Z(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n832), .B2(new_n833), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n827), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT102), .ZN(G145));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n507), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT103), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n496), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n691), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n746), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n758), .B(KEYINPUT104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n483), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n463), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n476), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(new_n797), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n623), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(G160), .B(new_n633), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n487), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n847), .A2(new_n854), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n847), .A2(KEYINPUT105), .A3(new_n854), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n857), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT106), .B1(new_n866), .B2(new_n857), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g447(.A(new_n830), .B(new_n616), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n604), .B(G299), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT107), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n876), .B1(new_n882), .B2(new_n873), .ZN(new_n883));
  XOR2_X1   g458(.A(G288), .B(G290), .Z(new_n884));
  XNOR2_X1  g459(.A(G305), .B(G303), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT42), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(KEYINPUT108), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n888), .B2(KEYINPUT42), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n883), .B(new_n889), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G868), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n824), .A2(new_n605), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  NAND2_X1  g468(.A1(G295), .A2(KEYINPUT109), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G331));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  XNOR2_X1  g473(.A(G301), .B(G286), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(new_n831), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n831), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(KEYINPUT110), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n901), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n906), .B2(new_n882), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n898), .B1(new_n907), .B2(new_n888), .ZN(new_n908));
  INV_X1    g483(.A(new_n888), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n903), .ZN(new_n910));
  INV_X1    g485(.A(new_n880), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n877), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n903), .B(new_n915), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n912), .A2(new_n913), .B1(new_n902), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n909), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n908), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n900), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n921), .A2(new_n881), .B1(new_n903), .B2(new_n902), .ZN(new_n922));
  AOI21_X1  g497(.A(G37), .B1(new_n922), .B2(new_n909), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n907), .A2(new_n888), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n908), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(KEYINPUT43), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n929), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g505(.A(KEYINPUT127), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n758), .B(new_n762), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n691), .B(G1996), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n797), .B(new_n799), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n843), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(G160), .A2(G40), .ZN(new_n945));
  OR3_X1    g520(.A1(new_n944), .A2(KEYINPUT112), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT112), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(G2078), .ZN(new_n954));
  INV_X1    g529(.A(G40), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n475), .A2(new_n480), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT124), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n509), .A2(new_n941), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n943), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(new_n443), .A3(new_n956), .A4(new_n951), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n952), .A2(new_n959), .B1(new_n962), .B2(new_n953), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n843), .A2(new_n964), .A3(new_n941), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n945), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n843), .A2(new_n968), .A3(new_n964), .A4(new_n941), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT123), .ZN(new_n971));
  INV_X1    g546(.A(G1961), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  OAI211_X1 g549(.A(G301), .B(new_n963), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n962), .A2(new_n953), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT122), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n496), .B2(new_n508), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n956), .B1(new_n979), .B2(new_n964), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(KEYINPUT114), .B2(new_n965), .ZN(new_n981));
  AOI21_X1  g556(.A(G1961), .B1(new_n981), .B2(new_n969), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n944), .A2(new_n956), .A3(new_n954), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n978), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n970), .A2(new_n972), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT122), .A3(new_n984), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n977), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n975), .B1(new_n989), .B2(G301), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT125), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n990), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n963), .B1(new_n973), .B2(new_n974), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n995), .B2(G171), .ZN(new_n996));
  INV_X1    g571(.A(new_n988), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT122), .B1(new_n987), .B2(new_n984), .ZN(new_n998));
  OAI211_X1 g573(.A(G301), .B(new_n976), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1981), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n580), .C1(new_n589), .C2(new_n593), .ZN(new_n1002));
  OAI21_X1  g577(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n580), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G1981), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(KEYINPUT49), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT115), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1002), .A2(new_n1011), .A3(KEYINPUT49), .A4(new_n1005), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  INV_X1    g588(.A(new_n842), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT103), .B1(new_n505), .B2(new_n506), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1016), .B2(new_n496), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1013), .B1(new_n1017), .B2(new_n956), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1007), .A2(new_n1010), .A3(new_n1012), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1018), .B(new_n1021), .C1(new_n1020), .C2(G288), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n843), .A2(new_n941), .A3(new_n956), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(G8), .C1(new_n1020), .C2(G288), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  NOR3_X1   g602(.A1(G166), .A2(new_n1027), .A3(new_n1013), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n961), .A2(new_n956), .A3(new_n951), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n781), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n966), .A2(new_n967), .A3(new_n1033), .A4(new_n969), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1026), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n945), .B1(new_n942), .B2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n979), .A2(KEYINPUT116), .A3(new_n964), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1038), .A2(new_n1033), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(new_n1032), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT117), .B(new_n1037), .C1(new_n1043), .C2(new_n1013), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1013), .B1(new_n1042), .B2(new_n1032), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1037), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1036), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n944), .A2(new_n956), .A3(new_n983), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n705), .ZN(new_n1051));
  INV_X1    g626(.A(G2084), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n966), .A2(new_n967), .A3(new_n1052), .A4(new_n969), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(G168), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(G168), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1058), .A3(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1000), .A2(new_n1049), .A3(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n993), .A2(new_n994), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1038), .A2(new_n1041), .A3(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT56), .B(G2072), .Z(new_n1066));
  OR2_X1    g641(.A1(new_n1031), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(G299), .B(KEYINPUT57), .Z(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1023), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1031), .B2(G1996), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n557), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT59), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT61), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1017), .A2(new_n1083), .A3(new_n762), .A4(new_n956), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n956), .A3(new_n941), .A4(new_n762), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1086));
  AOI221_X4 g661(.A(new_n1082), .B1(new_n1084), .B2(new_n1086), .C1(new_n970), .C2(new_n710), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n970), .A2(new_n710), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT121), .B(KEYINPUT60), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n612), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1348), .B1(new_n981), .B2(new_n969), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1082), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(KEYINPUT119), .A3(new_n1089), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT121), .B1(new_n1097), .B2(KEYINPUT60), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(new_n604), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1087), .A2(new_n1090), .A3(KEYINPUT60), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1081), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1095), .A2(new_n612), .A3(new_n1096), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1071), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n1072), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1072), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1109), .B(new_n1110), .C1(new_n1106), .C2(new_n1071), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1105), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1062), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n989), .A2(G301), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1057), .A2(new_n1117), .A3(new_n1059), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1049), .A4(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G168), .A2(G8), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(KEYINPUT63), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1049), .A2(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1026), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1037), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT63), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1030), .B(new_n1026), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1019), .A2(new_n1020), .A3(new_n577), .A4(new_n578), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1002), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1018), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1119), .A2(new_n1123), .A3(new_n1127), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n950), .B1(new_n1114), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n758), .A2(G2067), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n797), .A2(new_n800), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n934), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n949), .A2(new_n1137), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT48), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n948), .B2(new_n936), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n949), .B2(G1996), .ZN(new_n1146));
  INV_X1    g721(.A(G1996), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n948), .A2(KEYINPUT46), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n932), .A2(new_n691), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n948), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n931), .B1(new_n1134), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1155), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1132), .B1(new_n1113), .B2(new_n1062), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1157), .B(KEYINPUT127), .C1(new_n1158), .C2(new_n950), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1156), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g735(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n1162));
  OR2_X1    g736(.A1(new_n908), .A2(new_n918), .ZN(new_n1163));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1163), .B2(KEYINPUT43), .ZN(new_n1164));
  INV_X1    g738(.A(G319), .ZN(new_n1165));
  NOR4_X1   g739(.A1(G229), .A2(new_n1165), .A3(G401), .A4(G227), .ZN(new_n1166));
  AND3_X1   g740(.A1(new_n1164), .A2(new_n871), .A3(new_n1166), .ZN(G308));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n871), .A3(new_n1166), .ZN(G225));
endmodule


