

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760;

  OR2_X1 U372 ( .A1(n597), .A2(n624), .ZN(n450) );
  NAND2_X1 U373 ( .A1(n629), .A2(n628), .ZN(n624) );
  OR2_X1 U374 ( .A1(n709), .A2(G902), .ZN(n430) );
  XNOR2_X1 U375 ( .A(n491), .B(n490), .ZN(n498) );
  INV_X2 U376 ( .A(G146), .ZN(n434) );
  NAND2_X1 U377 ( .A1(n350), .A2(n360), .ZN(n395) );
  NAND2_X1 U378 ( .A1(n418), .A2(n417), .ZN(n350) );
  XNOR2_X1 U379 ( .A(n503), .B(n502), .ZN(n734) );
  NOR2_X2 U380 ( .A1(n703), .A2(n591), .ZN(n417) );
  NOR2_X2 U381 ( .A1(n607), .A2(n532), .ZN(n534) );
  OR2_X2 U382 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X2 U383 ( .A(G122), .B(G107), .ZN(n491) );
  NOR2_X2 U384 ( .A1(n583), .A2(n655), .ZN(n562) );
  NAND2_X1 U385 ( .A1(n367), .A2(n368), .ZN(n370) );
  NAND2_X1 U386 ( .A1(n738), .A2(n621), .ZN(n666) );
  NAND2_X1 U387 ( .A1(n402), .A2(n406), .ZN(n401) );
  AND2_X1 U388 ( .A1(n400), .A2(n399), .ZN(n398) );
  OR2_X1 U389 ( .A1(n635), .A2(n576), .ZN(n577) );
  XOR2_X1 U390 ( .A(KEYINPUT62), .B(n680), .Z(n681) );
  XNOR2_X1 U391 ( .A(n374), .B(n373), .ZN(n486) );
  XNOR2_X1 U392 ( .A(n416), .B(G137), .ZN(n431) );
  NAND2_X1 U393 ( .A1(n393), .A2(n392), .ZN(n351) );
  NAND2_X1 U394 ( .A1(n393), .A2(n392), .ZN(n396) );
  XNOR2_X1 U395 ( .A(n372), .B(n363), .ZN(n615) );
  NAND2_X1 U396 ( .A1(n615), .A2(n614), .ZN(n620) );
  NOR2_X1 U397 ( .A1(n607), .A2(n532), .ZN(n352) );
  NOR2_X1 U398 ( .A1(n671), .A2(n670), .ZN(n353) );
  XNOR2_X1 U399 ( .A(n396), .B(n364), .ZN(n354) );
  NOR2_X1 U400 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U401 ( .A(n351), .B(n364), .ZN(n667) );
  XNOR2_X1 U402 ( .A(n550), .B(KEYINPUT109), .ZN(n603) );
  NOR2_X1 U403 ( .A1(G953), .A2(G237), .ZN(n471) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n514) );
  NOR2_X1 U405 ( .A1(n663), .A2(n390), .ZN(n389) );
  NAND2_X1 U406 ( .A1(n610), .A2(n391), .ZN(n390) );
  XNOR2_X1 U407 ( .A(n519), .B(KEYINPUT38), .ZN(n593) );
  NAND2_X1 U408 ( .A1(n515), .A2(G214), .ZN(n641) );
  XNOR2_X1 U409 ( .A(n469), .B(KEYINPUT81), .ZN(n544) );
  XNOR2_X1 U410 ( .A(n497), .B(n496), .ZN(n535) );
  XNOR2_X1 U411 ( .A(n485), .B(n484), .ZN(n536) );
  XNOR2_X1 U412 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U413 ( .A(KEYINPUT0), .ZN(n533) );
  INV_X2 U414 ( .A(G953), .ZN(n752) );
  XNOR2_X1 U415 ( .A(n498), .B(n376), .ZN(n503) );
  XNOR2_X1 U416 ( .A(n603), .B(n602), .ZN(n415) );
  NAND2_X1 U417 ( .A1(n412), .A2(KEYINPUT36), .ZN(n411) );
  NAND2_X1 U418 ( .A1(n387), .A2(n388), .ZN(n386) );
  INV_X1 U419 ( .A(KEYINPUT46), .ZN(n385) );
  XNOR2_X1 U420 ( .A(KEYINPUT72), .B(G131), .ZN(n478) );
  AND2_X1 U421 ( .A1(n355), .A2(n588), .ZN(n375) );
  XNOR2_X1 U422 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n452) );
  INV_X1 U423 ( .A(G137), .ZN(n451) );
  XNOR2_X1 U424 ( .A(KEYINPUT3), .B(G119), .ZN(n499) );
  XNOR2_X1 U425 ( .A(G113), .B(G116), .ZN(n456) );
  INV_X1 U426 ( .A(n499), .ZN(n376) );
  XNOR2_X1 U427 ( .A(G104), .B(G113), .ZN(n501) );
  XOR2_X1 U428 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n473) );
  XNOR2_X1 U429 ( .A(G140), .B(G143), .ZN(n474) );
  XOR2_X1 U430 ( .A(KEYINPUT12), .B(G122), .Z(n475) );
  INV_X1 U431 ( .A(G140), .ZN(n416) );
  XOR2_X1 U432 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n510) );
  XNOR2_X1 U433 ( .A(n383), .B(n361), .ZN(n466) );
  XNOR2_X1 U434 ( .A(KEYINPUT14), .B(KEYINPUT91), .ZN(n383) );
  NOR2_X1 U435 ( .A1(n593), .A2(n544), .ZN(n405) );
  INV_X1 U436 ( .A(KEYINPUT39), .ZN(n407) );
  NAND2_X1 U437 ( .A1(n470), .A2(n407), .ZN(n399) );
  XOR2_X1 U438 ( .A(n516), .B(KEYINPUT90), .Z(n517) );
  INV_X1 U439 ( .A(G902), .ZN(n495) );
  INV_X1 U440 ( .A(KEYINPUT8), .ZN(n373) );
  NAND2_X1 U441 ( .A1(n752), .A2(G234), .ZN(n374) );
  INV_X1 U442 ( .A(G116), .ZN(n490) );
  BUF_X1 U443 ( .A(n668), .Z(n751) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n420) );
  INV_X1 U445 ( .A(KEYINPUT92), .ZN(n381) );
  NAND2_X1 U446 ( .A1(n466), .A2(G952), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n560), .B(n559), .ZN(n655) );
  XNOR2_X1 U448 ( .A(n594), .B(KEYINPUT41), .ZN(n656) );
  XNOR2_X1 U449 ( .A(n378), .B(KEYINPUT74), .ZN(n595) );
  NAND2_X1 U450 ( .A1(n380), .A2(n359), .ZN(n378) );
  INV_X1 U451 ( .A(n544), .ZN(n403) );
  INV_X1 U452 ( .A(n470), .ZN(n406) );
  XNOR2_X1 U453 ( .A(n538), .B(KEYINPUT22), .ZN(n571) );
  XNOR2_X1 U454 ( .A(n634), .B(KEYINPUT6), .ZN(n567) );
  XNOR2_X1 U455 ( .A(n687), .B(n686), .ZN(n688) );
  INV_X1 U456 ( .A(KEYINPUT64), .ZN(n368) );
  XNOR2_X1 U457 ( .A(n696), .B(n695), .ZN(n697) );
  AND2_X1 U458 ( .A1(n411), .A2(n558), .ZN(n410) );
  AND2_X1 U459 ( .A1(n704), .A2(n573), .ZN(n355) );
  AND2_X1 U460 ( .A1(n573), .A2(n397), .ZN(n356) );
  INV_X1 U461 ( .A(n628), .ZN(n379) );
  OR2_X1 U462 ( .A1(G902), .A2(G237), .ZN(n357) );
  XOR2_X1 U463 ( .A(n489), .B(KEYINPUT9), .Z(n358) );
  NOR2_X1 U464 ( .A1(n544), .A2(n379), .ZN(n359) );
  OR2_X1 U465 ( .A1(n591), .A2(n590), .ZN(n360) );
  AND2_X1 U466 ( .A1(G234), .A2(G237), .ZN(n361) );
  AND2_X1 U467 ( .A1(n581), .A2(n403), .ZN(n362) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n414) );
  XOR2_X1 U469 ( .A(n611), .B(KEYINPUT73), .Z(n363) );
  XNOR2_X1 U470 ( .A(KEYINPUT87), .B(KEYINPUT45), .ZN(n364) );
  XNOR2_X1 U471 ( .A(n352), .B(n533), .ZN(n365) );
  XNOR2_X1 U472 ( .A(n565), .B(KEYINPUT35), .ZN(n366) );
  NAND2_X1 U473 ( .A1(n353), .A2(KEYINPUT64), .ZN(n369) );
  NAND2_X2 U474 ( .A1(n370), .A2(n369), .ZN(n705) );
  INV_X1 U475 ( .A(n672), .ZN(n367) );
  XNOR2_X1 U476 ( .A(n534), .B(n533), .ZN(n578) );
  XNOR2_X1 U477 ( .A(n565), .B(KEYINPUT35), .ZN(n703) );
  XNOR2_X1 U478 ( .A(n423), .B(G146), .ZN(n455) );
  INV_X1 U479 ( .A(n605), .ZN(n412) );
  OR2_X1 U480 ( .A1(n365), .A2(n577), .ZN(n580) );
  NAND2_X1 U481 ( .A1(n575), .A2(n574), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n386), .B(n385), .ZN(n384) );
  NAND2_X1 U483 ( .A1(n384), .A2(n389), .ZN(n372) );
  XNOR2_X1 U484 ( .A(n432), .B(n433), .ZN(n440) );
  XNOR2_X1 U485 ( .A(n620), .B(KEYINPUT86), .ZN(n668) );
  NAND2_X1 U486 ( .A1(n566), .A2(n375), .ZN(n392) );
  XNOR2_X1 U487 ( .A(n513), .B(n734), .ZN(n693) );
  NAND2_X1 U488 ( .A1(n377), .A2(n410), .ZN(n409) );
  NAND2_X1 U489 ( .A1(n415), .A2(n413), .ZN(n377) );
  INV_X1 U490 ( .A(n629), .ZN(n380) );
  XNOR2_X2 U491 ( .A(n447), .B(n446), .ZN(n629) );
  INV_X1 U492 ( .A(n601), .ZN(n387) );
  INV_X1 U493 ( .A(n760), .ZN(n388) );
  INV_X1 U494 ( .A(n606), .ZN(n391) );
  NAND2_X1 U495 ( .A1(n355), .A2(KEYINPUT65), .ZN(n394) );
  AND2_X2 U496 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U497 ( .A1(n704), .A2(n356), .ZN(n575) );
  INV_X1 U498 ( .A(KEYINPUT69), .ZN(n397) );
  XNOR2_X2 U499 ( .A(n572), .B(KEYINPUT32), .ZN(n704) );
  NAND2_X1 U500 ( .A1(n401), .A2(n398), .ZN(n555) );
  NAND2_X1 U501 ( .A1(n404), .A2(n407), .ZN(n400) );
  NOR2_X1 U502 ( .A1(n404), .A2(n407), .ZN(n402) );
  NAND2_X1 U503 ( .A1(n406), .A2(n362), .ZN(n521) );
  NAND2_X1 U504 ( .A1(n581), .A2(n405), .ZN(n404) );
  XNOR2_X2 U505 ( .A(n450), .B(KEYINPUT99), .ZN(n581) );
  NOR2_X1 U506 ( .A1(n409), .A2(n408), .ZN(n663) );
  NOR2_X1 U507 ( .A1(n415), .A2(n414), .ZN(n408) );
  AND2_X1 U508 ( .A1(n605), .A2(n414), .ZN(n413) );
  XNOR2_X2 U509 ( .A(KEYINPUT68), .B(G101), .ZN(n423) );
  INV_X1 U510 ( .A(n634), .ZN(n576) );
  NAND2_X1 U511 ( .A1(n634), .A2(n641), .ZN(n465) );
  XNOR2_X2 U512 ( .A(n463), .B(G472), .ZN(n634) );
  NOR2_X2 U513 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X2 U514 ( .A1(n525), .A2(n641), .ZN(n526) );
  XNOR2_X2 U515 ( .A(n518), .B(n517), .ZN(n525) );
  NAND2_X1 U516 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U517 ( .A1(n643), .A2(n379), .ZN(n419) );
  INV_X1 U518 ( .A(KEYINPUT111), .ZN(n602) );
  XNOR2_X2 U519 ( .A(G143), .B(G128), .ZN(n492) );
  XNOR2_X1 U520 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n421) );
  XNOR2_X1 U521 ( .A(n492), .B(n421), .ZN(n506) );
  XNOR2_X1 U522 ( .A(n478), .B(G134), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n506), .B(n422), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n461), .B(n431), .ZN(n750) );
  NAND2_X1 U525 ( .A1(n752), .A2(G227), .ZN(n424) );
  XNOR2_X1 U526 ( .A(n424), .B(G110), .ZN(n426) );
  XNOR2_X1 U527 ( .A(G104), .B(G107), .ZN(n425) );
  XNOR2_X1 U528 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n455), .B(n427), .ZN(n428) );
  XNOR2_X1 U530 ( .A(n750), .B(n428), .ZN(n709) );
  XNOR2_X1 U531 ( .A(KEYINPUT75), .B(G469), .ZN(n429) );
  XNOR2_X2 U532 ( .A(n430), .B(n429), .ZN(n597) );
  XOR2_X1 U533 ( .A(n431), .B(KEYINPUT24), .Z(n433) );
  NAND2_X1 U534 ( .A1(G221), .A2(n486), .ZN(n432) );
  XNOR2_X2 U535 ( .A(n434), .B(G125), .ZN(n505) );
  XNOR2_X1 U536 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U537 ( .A(n505), .B(n435), .ZN(n749) );
  XOR2_X1 U538 ( .A(KEYINPUT23), .B(G119), .Z(n437) );
  XNOR2_X1 U539 ( .A(G128), .B(G110), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n438), .B(n749), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n440), .B(n439), .ZN(n678) );
  NAND2_X1 U543 ( .A1(n678), .A2(n495), .ZN(n447) );
  XNOR2_X1 U544 ( .A(KEYINPUT78), .B(KEYINPUT97), .ZN(n443) );
  NAND2_X1 U545 ( .A1(G234), .A2(n514), .ZN(n441) );
  XNOR2_X1 U546 ( .A(KEYINPUT20), .B(n441), .ZN(n448) );
  AND2_X1 U547 ( .A1(n448), .A2(G217), .ZN(n442) );
  XNOR2_X1 U548 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U549 ( .A(KEYINPUT25), .B(KEYINPUT98), .Z(n444) );
  XNOR2_X1 U550 ( .A(n445), .B(n444), .ZN(n446) );
  AND2_X1 U551 ( .A1(n448), .A2(G221), .ZN(n449) );
  XNOR2_X1 U552 ( .A(n449), .B(KEYINPUT21), .ZN(n628) );
  XNOR2_X1 U553 ( .A(n451), .B(KEYINPUT100), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U555 ( .A(n455), .B(n454), .ZN(n460) );
  NAND2_X1 U556 ( .A1(n471), .A2(G210), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U558 ( .A(n458), .B(n499), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U560 ( .A(n461), .B(n462), .ZN(n680) );
  OR2_X1 U561 ( .A1(n680), .A2(G902), .ZN(n463) );
  XNOR2_X1 U562 ( .A(KEYINPUT76), .B(n357), .ZN(n515) );
  XNOR2_X1 U563 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n464) );
  XNOR2_X1 U564 ( .A(n465), .B(n464), .ZN(n470) );
  NAND2_X1 U565 ( .A1(n420), .A2(n752), .ZN(n531) );
  NAND2_X1 U566 ( .A1(G902), .A2(n466), .ZN(n528) );
  NOR2_X1 U567 ( .A1(G900), .A2(n528), .ZN(n467) );
  NAND2_X1 U568 ( .A1(n467), .A2(G953), .ZN(n468) );
  NAND2_X1 U569 ( .A1(n531), .A2(n468), .ZN(n469) );
  NAND2_X1 U570 ( .A1(n471), .A2(G214), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U573 ( .A(n477), .B(n476), .Z(n481) );
  XOR2_X1 U574 ( .A(n478), .B(n501), .Z(n479) );
  XNOR2_X1 U575 ( .A(n749), .B(n479), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n481), .B(n480), .ZN(n687) );
  NOR2_X1 U577 ( .A1(G902), .A2(n687), .ZN(n485) );
  XNOR2_X1 U578 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n483) );
  INV_X1 U579 ( .A(G475), .ZN(n482) );
  XOR2_X1 U580 ( .A(G134), .B(KEYINPUT104), .Z(n488) );
  NAND2_X1 U581 ( .A1(G217), .A2(n486), .ZN(n487) );
  XNOR2_X1 U582 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n492), .B(KEYINPUT7), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n498), .B(n493), .ZN(n494) );
  XNOR2_X1 U585 ( .A(n358), .B(n494), .ZN(n674) );
  NAND2_X1 U586 ( .A1(n674), .A2(n495), .ZN(n497) );
  XNOR2_X1 U587 ( .A(KEYINPUT105), .B(G478), .ZN(n496) );
  NOR2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n563) );
  XNOR2_X1 U589 ( .A(G110), .B(KEYINPUT16), .ZN(n500) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U591 ( .A(n423), .ZN(n504) );
  XNOR2_X1 U592 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n507), .B(n506), .ZN(n512) );
  NAND2_X1 U594 ( .A1(G224), .A2(n752), .ZN(n508) );
  XNOR2_X1 U595 ( .A(n508), .B(KEYINPUT79), .ZN(n509) );
  XNOR2_X1 U596 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U597 ( .A(n512), .B(n511), .ZN(n513) );
  INV_X1 U598 ( .A(n514), .ZN(n665) );
  NOR2_X2 U599 ( .A1(n693), .A2(n665), .ZN(n518) );
  AND2_X1 U600 ( .A1(n515), .A2(G210), .ZN(n516) );
  BUF_X1 U601 ( .A(n525), .Z(n519) );
  NAND2_X1 U602 ( .A1(n563), .A2(n519), .ZN(n520) );
  NOR2_X1 U603 ( .A1(n521), .A2(n520), .ZN(n606) );
  XOR2_X1 U604 ( .A(G143), .B(n606), .Z(G45) );
  INV_X1 U605 ( .A(KEYINPUT103), .ZN(n522) );
  XNOR2_X1 U606 ( .A(n536), .B(n522), .ZN(n547) );
  INV_X1 U607 ( .A(n535), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n524) );
  INV_X1 U609 ( .A(KEYINPUT107), .ZN(n523) );
  XNOR2_X1 U610 ( .A(n524), .B(n523), .ZN(n732) );
  NOR2_X1 U611 ( .A1(n555), .A2(n732), .ZN(n612) );
  XOR2_X1 U612 ( .A(G134), .B(n612), .Z(G36) );
  XNOR2_X2 U613 ( .A(n526), .B(KEYINPUT89), .ZN(n604) );
  XNOR2_X2 U614 ( .A(n604), .B(KEYINPUT19), .ZN(n607) );
  XNOR2_X1 U615 ( .A(G898), .B(KEYINPUT93), .ZN(n743) );
  NAND2_X1 U616 ( .A1(n743), .A2(G953), .ZN(n527) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT94), .ZN(n736) );
  NOR2_X1 U618 ( .A1(n736), .A2(n528), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n529), .B(KEYINPUT95), .ZN(n530) );
  AND2_X1 U620 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U621 ( .A(n365), .ZN(n537) );
  NAND2_X1 U622 ( .A1(n536), .A2(n535), .ZN(n643) );
  NAND2_X1 U623 ( .A1(n537), .A2(n419), .ZN(n538) );
  XNOR2_X2 U624 ( .A(n597), .B(KEYINPUT1), .ZN(n625) );
  NOR2_X1 U625 ( .A1(n634), .A2(n629), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n625), .A2(n539), .ZN(n540) );
  OR2_X1 U627 ( .A1(n571), .A2(n540), .ZN(n573) );
  XOR2_X1 U628 ( .A(G110), .B(KEYINPUT113), .Z(n541) );
  XNOR2_X1 U629 ( .A(n573), .B(n541), .ZN(G12) );
  AND2_X1 U630 ( .A1(n567), .A2(n629), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n625), .A2(n542), .ZN(n543) );
  OR2_X1 U632 ( .A1(n571), .A2(n543), .ZN(n586) );
  XNOR2_X1 U633 ( .A(n586), .B(G101), .ZN(G3) );
  NOR2_X1 U634 ( .A1(n595), .A2(n567), .ZN(n545) );
  XNOR2_X1 U635 ( .A(KEYINPUT108), .B(n545), .ZN(n549) );
  NOR2_X1 U636 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n548), .B(KEYINPUT106), .ZN(n724) );
  NAND2_X1 U638 ( .A1(n549), .A2(n724), .ZN(n550) );
  INV_X1 U639 ( .A(n625), .ZN(n558) );
  INV_X1 U640 ( .A(n641), .ZN(n551) );
  NOR2_X1 U641 ( .A1(n558), .A2(n551), .ZN(n552) );
  NAND2_X1 U642 ( .A1(n603), .A2(n552), .ZN(n553) );
  XOR2_X1 U643 ( .A(KEYINPUT43), .B(n553), .Z(n554) );
  NOR2_X1 U644 ( .A1(n554), .A2(n519), .ZN(n613) );
  XOR2_X1 U645 ( .A(G140), .B(n613), .Z(G42) );
  INV_X1 U646 ( .A(n724), .ZN(n728) );
  NOR2_X1 U647 ( .A1(n555), .A2(n728), .ZN(n556) );
  XNOR2_X1 U648 ( .A(n556), .B(KEYINPUT40), .ZN(n601) );
  XOR2_X1 U649 ( .A(n601), .B(G131), .Z(G33) );
  XNOR2_X1 U650 ( .A(n578), .B(KEYINPUT96), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n624), .A2(n567), .ZN(n557) );
  NAND2_X1 U652 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U653 ( .A(KEYINPUT33), .ZN(n559) );
  XNOR2_X1 U654 ( .A(KEYINPUT80), .B(KEYINPUT34), .ZN(n561) );
  XNOR2_X1 U655 ( .A(n562), .B(n561), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n366), .B(KEYINPUT69), .ZN(n566) );
  INV_X1 U657 ( .A(KEYINPUT44), .ZN(n588) );
  INV_X1 U658 ( .A(n567), .ZN(n568) );
  OR2_X1 U659 ( .A1(n568), .A2(n629), .ZN(n569) );
  OR2_X1 U660 ( .A1(n625), .A2(n569), .ZN(n570) );
  INV_X1 U661 ( .A(KEYINPUT65), .ZN(n589) );
  OR2_X1 U662 ( .A1(n588), .A2(n589), .ZN(n574) );
  OR2_X1 U663 ( .A1(n625), .A2(n624), .ZN(n635) );
  INV_X1 U664 ( .A(KEYINPUT31), .ZN(n579) );
  XNOR2_X2 U665 ( .A(n580), .B(n579), .ZN(n731) );
  NAND2_X1 U666 ( .A1(n581), .A2(n576), .ZN(n582) );
  OR2_X1 U667 ( .A1(n583), .A2(n582), .ZN(n717) );
  NAND2_X1 U668 ( .A1(n731), .A2(n717), .ZN(n585) );
  AND2_X1 U669 ( .A1(n732), .A2(n728), .ZN(n647) );
  INV_X1 U670 ( .A(n647), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U672 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U674 ( .A(KEYINPUT2), .ZN(n619) );
  NAND2_X1 U675 ( .A1(n354), .A2(n619), .ZN(n592) );
  XNOR2_X1 U676 ( .A(n592), .B(KEYINPUT84), .ZN(n617) );
  INV_X1 U677 ( .A(n593), .ZN(n642) );
  NAND2_X1 U678 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U679 ( .A1(n643), .A2(n646), .ZN(n594) );
  NOR2_X1 U680 ( .A1(n595), .A2(n576), .ZN(n596) );
  XNOR2_X1 U681 ( .A(n596), .B(KEYINPUT28), .ZN(n599) );
  INV_X1 U682 ( .A(n597), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n723) );
  NOR2_X1 U684 ( .A1(n656), .A2(n723), .ZN(n600) );
  XNOR2_X1 U685 ( .A(n600), .B(KEYINPUT42), .ZN(n760) );
  BUF_X1 U686 ( .A(n604), .Z(n605) );
  BUF_X1 U687 ( .A(n607), .Z(n608) );
  OR2_X1 U688 ( .A1(n723), .A2(n608), .ZN(n720) );
  NOR2_X1 U689 ( .A1(n720), .A2(n647), .ZN(n609) );
  XNOR2_X1 U690 ( .A(n609), .B(KEYINPUT47), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n611) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n751), .A2(n619), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT82), .B(n618), .Z(n622) );
  INV_X1 U696 ( .A(n667), .ZN(n738) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n666), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT85), .ZN(n661) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  XOR2_X1 U701 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n626) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(n632) );
  NOR2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(KEYINPUT49), .B(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U706 ( .A1(n633), .A2(n576), .ZN(n637) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT51), .B(n638), .Z(n639) );
  NOR2_X1 U710 ( .A1(n656), .A2(n639), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n640), .B(KEYINPUT116), .ZN(n652) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U714 ( .A(KEYINPUT117), .B(n645), .Z(n649) );
  NOR2_X1 U715 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n650), .A2(n655), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U719 ( .A(KEYINPUT52), .B(n653), .Z(n654) );
  NAND2_X1 U720 ( .A1(n654), .A2(n420), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n657), .A2(G953), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U724 ( .A(n662), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U725 ( .A(G125), .B(KEYINPUT37), .Z(n664) );
  XOR2_X1 U726 ( .A(n664), .B(n663), .Z(G27) );
  NAND2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n671) );
  NOR2_X1 U728 ( .A1(n668), .A2(n354), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n669), .A2(KEYINPUT2), .ZN(n670) );
  NAND2_X1 U730 ( .A1(n705), .A2(G478), .ZN(n673) );
  XOR2_X1 U731 ( .A(n674), .B(n673), .Z(n676) );
  INV_X1 U732 ( .A(G952), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n675), .A2(G953), .ZN(n699) );
  INV_X1 U734 ( .A(n699), .ZN(n712) );
  NOR2_X1 U735 ( .A1(n676), .A2(n712), .ZN(G63) );
  NAND2_X1 U736 ( .A1(n705), .A2(G217), .ZN(n677) );
  XOR2_X1 U737 ( .A(n678), .B(n677), .Z(n679) );
  NOR2_X1 U738 ( .A1(n679), .A2(n712), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n705), .A2(G472), .ZN(n682) );
  XNOR2_X1 U740 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U741 ( .A1(n683), .A2(n699), .ZN(n684) );
  XNOR2_X1 U742 ( .A(n684), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U743 ( .A1(n705), .A2(G475), .ZN(n689) );
  XNOR2_X1 U744 ( .A(KEYINPUT66), .B(KEYINPUT121), .ZN(n685) );
  XOR2_X1 U745 ( .A(n685), .B(KEYINPUT59), .Z(n686) );
  XNOR2_X1 U746 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U747 ( .A1(n690), .A2(n699), .ZN(n692) );
  XNOR2_X1 U748 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n692), .B(n691), .ZN(G60) );
  NAND2_X1 U750 ( .A1(n705), .A2(G210), .ZN(n698) );
  BUF_X1 U751 ( .A(n693), .Z(n696) );
  XNOR2_X1 U752 ( .A(KEYINPUT83), .B(KEYINPUT54), .ZN(n694) );
  XOR2_X1 U753 ( .A(n694), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U756 ( .A(KEYINPUT118), .B(KEYINPUT56), .Z(n701) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(G51) );
  XOR2_X1 U758 ( .A(n366), .B(G122), .Z(G24) );
  XNOR2_X1 U759 ( .A(n704), .B(G119), .ZN(G21) );
  NAND2_X1 U760 ( .A1(n705), .A2(G469), .ZN(n711) );
  XNOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n707) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n706) );
  XNOR2_X1 U763 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(G54) );
  NOR2_X1 U767 ( .A1(n717), .A2(n728), .ZN(n714) );
  XOR2_X1 U768 ( .A(G104), .B(n714), .Z(G6) );
  XOR2_X1 U769 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n716) );
  XNOR2_X1 U770 ( .A(G107), .B(KEYINPUT27), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n719) );
  NOR2_X1 U772 ( .A1(n717), .A2(n732), .ZN(n718) );
  XOR2_X1 U773 ( .A(n719), .B(n718), .Z(G9) );
  NOR2_X1 U774 ( .A1(n720), .A2(n732), .ZN(n722) );
  XNOR2_X1 U775 ( .A(G128), .B(KEYINPUT29), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n722), .B(n721), .ZN(G30) );
  INV_X1 U777 ( .A(n723), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n726), .A2(n608), .ZN(n727) );
  XOR2_X1 U780 ( .A(G146), .B(n727), .Z(G48) );
  NOR2_X1 U781 ( .A1(n728), .A2(n731), .ZN(n729) );
  XOR2_X1 U782 ( .A(KEYINPUT114), .B(n729), .Z(n730) );
  XNOR2_X1 U783 ( .A(G113), .B(n730), .ZN(G15) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U785 ( .A(G116), .B(n733), .Z(G18) );
  XNOR2_X1 U786 ( .A(G101), .B(KEYINPUT125), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n734), .B(n735), .ZN(n737) );
  NAND2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n747) );
  NAND2_X1 U789 ( .A1(n738), .A2(n752), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(KEYINPUT123), .ZN(n745) );
  XOR2_X1 U791 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n741) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n740) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U795 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U797 ( .A(KEYINPUT124), .B(n748), .ZN(G69) );
  XNOR2_X1 U798 ( .A(n750), .B(n749), .ZN(n755) );
  XNOR2_X1 U799 ( .A(n751), .B(n755), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT126), .ZN(n759) );
  XNOR2_X1 U802 ( .A(n755), .B(G227), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(G72) );
  XOR2_X1 U806 ( .A(n760), .B(G137), .Z(G39) );
endmodule

