//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT11), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n187), .B(new_n192), .C1(new_n188), .C2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n196), .A3(new_n191), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(G104), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n200), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT76), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(new_n199), .A3(KEYINPUT76), .A4(G104), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT78), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n199), .B2(G104), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n199), .A3(G104), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(KEYINPUT79), .A3(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G146), .ZN(new_n225));
  AND4_X1   g039(.A1(new_n221), .A2(new_n223), .A3(new_n225), .A4(G128), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g043(.A(G143), .B(G146), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n224), .B2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n225), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n220), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(KEYINPUT80), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(new_n240), .A3(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(G128), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n226), .B1(new_n242), .B2(new_n235), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n219), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n198), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n201), .A2(new_n203), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n210), .A2(G107), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n208), .A3(new_n207), .A4(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n250), .B2(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(KEYINPUT77), .A3(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(KEYINPUT77), .A3(KEYINPUT4), .A4(G101), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n235), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n219), .B2(new_n243), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(KEYINPUT81), .B(new_n260), .C1(new_n219), .C2(new_n243), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n237), .ZN(new_n265));
  AND4_X1   g079(.A1(new_n259), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n198), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT82), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n259), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n269), .A2(new_n270), .A3(new_n198), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n247), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n267), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n270), .B1(new_n269), .B2(new_n198), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n198), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n276), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT83), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n276), .B(new_n247), .C1(new_n268), .C2(new_n271), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n279), .A2(new_n280), .B1(new_n198), .B2(new_n269), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n276), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT84), .A2(G469), .ZN(new_n291));
  OR2_X1    g105(.A1(KEYINPUT84), .A2(G469), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n289), .A2(new_n290), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n277), .A2(new_n272), .B1(new_n295), .B2(new_n282), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(G469), .C1(new_n296), .C2(G902), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n300));
  INV_X1    g114(.A(G113), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT68), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT2), .A3(G113), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n302), .A2(new_n304), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  XNOR2_X1  g119(.A(G116), .B(G119), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n309), .A2(KEYINPUT5), .A3(G119), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(G113), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n219), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n305), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n255), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(G110), .B(G122), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT85), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n299), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n320), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n316), .B1(new_n253), .B2(new_n254), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT6), .B(new_n321), .C1(new_n325), .C2(new_n313), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n258), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n237), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT86), .B(G224), .Z(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n274), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n333), .A3(new_n330), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n327), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n335), .B(new_n336), .C1(KEYINPUT7), .C2(new_n334), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT88), .B1(new_n219), .B2(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n341), .A2(new_n312), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n341), .B(new_n312), .C1(KEYINPUT88), .C2(new_n219), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n319), .A2(KEYINPUT8), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n319), .A2(KEYINPUT8), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  OR3_X1    g160(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n334), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n339), .A2(new_n324), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G210), .B1(G237), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n338), .A2(new_n350), .A3(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(KEYINPUT89), .A3(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n353), .A2(KEYINPUT89), .ZN(new_n355));
  OAI21_X1  g169(.A(G214), .B1(G237), .B2(G902), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G221), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT9), .B(G234), .Z(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n290), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT75), .Z(new_n361));
  XNOR2_X1  g175(.A(G113), .B(G122), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(new_n210), .ZN(new_n363));
  NOR2_X1   g177(.A1(G237), .A2(G953), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G214), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT90), .A3(G143), .ZN(new_n366));
  OR2_X1    g180(.A1(KEYINPUT90), .A2(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT90), .A2(G143), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(G214), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT18), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n196), .ZN(new_n372));
  XNOR2_X1  g186(.A(G125), .B(G140), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n222), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n366), .A2(G131), .A3(new_n369), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n372), .B(new_n374), .C1(new_n371), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(G131), .B1(new_n366), .B2(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  INV_X1    g194(.A(new_n375), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n329), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(G146), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n222), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT72), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n384), .A2(new_n390), .A3(G146), .A4(new_n385), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n363), .B(new_n376), .C1(new_n383), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n373), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT19), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT19), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n373), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n222), .A3(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(new_n386), .C1(new_n381), .C2(new_n377), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n376), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n363), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G475), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n290), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT20), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n407), .A3(new_n404), .A4(new_n290), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n376), .B1(new_n383), .B2(new_n392), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n401), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n393), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n290), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G475), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G128), .B(G143), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT13), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n224), .A3(G128), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(G134), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n188), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(G107), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT91), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n199), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n420), .A4(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT14), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n309), .A2(KEYINPUT14), .A3(G122), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G107), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n423), .A2(new_n199), .ZN(new_n434));
  INV_X1    g248(.A(new_n421), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n416), .A2(new_n188), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n433), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n359), .A2(G217), .A3(new_n274), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n429), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n429), .B2(new_n437), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT92), .B(new_n290), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n188), .B1(new_n416), .B2(KEYINPUT13), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n435), .B1(new_n419), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n427), .B1(new_n447), .B2(new_n426), .ZN(new_n448));
  INV_X1    g262(.A(new_n428), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n437), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n438), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n429), .A2(new_n437), .A3(new_n439), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n444), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(KEYINPUT92), .A3(new_n290), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(G234), .A2(G237), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(G952), .A3(new_n274), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT21), .B(G898), .Z(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(G902), .A3(G953), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n415), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n298), .A2(new_n357), .A3(new_n361), .A4(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n191), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n188), .A2(G137), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n197), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n237), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT70), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n258), .A2(new_n198), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n237), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n317), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n470), .A2(new_n316), .A3(new_n471), .A4(new_n473), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT28), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n316), .A3(new_n469), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n364), .A2(G210), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT26), .B(G101), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(KEYINPUT30), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n197), .A2(KEYINPUT65), .A3(new_n467), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT65), .B1(new_n197), .B2(new_n467), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n237), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT67), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  OAI211_X1 g313(.A(KEYINPUT67), .B(new_n237), .C1(new_n494), .C2(new_n495), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n471), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n316), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n476), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n489), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n471), .A3(new_n500), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n503), .B1(new_n317), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n481), .B1(new_n506), .B2(new_n480), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n490), .B(new_n504), .C1(new_n507), .C2(new_n489), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n492), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G472), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  NOR2_X1   g325(.A1(G472), .A2(G902), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n317), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n480), .B1(new_n513), .B2(new_n476), .ZN(new_n514));
  INV_X1    g328(.A(new_n481), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n489), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n493), .A2(new_n501), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n317), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n476), .A4(new_n488), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n502), .A2(new_n503), .A3(new_n489), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n519), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n511), .B(new_n512), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n476), .A3(new_n488), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT31), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n520), .A3(new_n516), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n511), .B1(new_n528), .B2(new_n512), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n510), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G119), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G128), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(G128), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT24), .B(G110), .Z(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n534), .A2(KEYINPUT23), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(KEYINPUT23), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G110), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n392), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n540), .A2(G110), .B1(new_n535), .B2(new_n536), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n386), .C1(G146), .C2(new_n394), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n546), .B(new_n547), .Z(new_n548));
  XNOR2_X1  g362(.A(new_n545), .B(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n549), .A2(new_n290), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT25), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT74), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(KEYINPUT74), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G217), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(G234), .B2(new_n290), .ZN(new_n557));
  INV_X1    g371(.A(new_n553), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n555), .B(new_n557), .C1(new_n550), .C2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n549), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n530), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n464), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n205), .ZN(G3));
  NAND2_X1  g380(.A1(new_n528), .A2(new_n290), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n567), .A2(G472), .B1(new_n512), .B2(new_n528), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n298), .A2(new_n563), .A3(new_n361), .A4(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n338), .A2(new_n350), .A3(new_n348), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n350), .B1(new_n338), .B2(new_n348), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n356), .B(new_n461), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(new_n440), .B2(new_n441), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n453), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n443), .B(G902), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G478), .B1(new_n453), .B2(new_n290), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n415), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n571), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n356), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n352), .B2(new_n353), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n575), .A2(new_n576), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT33), .B1(new_n453), .B2(KEYINPUT93), .ZN(new_n586));
  OAI211_X1 g400(.A(G478), .B(new_n290), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n580), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n587), .A2(new_n588), .B1(new_n414), .B2(new_n409), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n584), .A2(KEYINPUT94), .A3(new_n461), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n570), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT34), .B(G104), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n411), .B2(new_n393), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n404), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n413), .A2(KEYINPUT95), .A3(G475), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n409), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n456), .A4(new_n461), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n409), .A2(new_n456), .A3(new_n598), .A4(new_n597), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT96), .B1(new_n602), .B2(new_n462), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n601), .A2(new_n603), .A3(new_n584), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n570), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(new_n199), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  INV_X1    g422(.A(new_n568), .ZN(new_n609));
  INV_X1    g423(.A(new_n548), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n545), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n560), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n559), .A2(new_n613), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n464), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT37), .B(G110), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G12));
  NAND2_X1  g431(.A1(new_n559), .A2(new_n613), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n618), .A2(new_n584), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n530), .A2(new_n298), .A3(new_n619), .A4(new_n361), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n458), .B1(new_n460), .B2(G900), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n602), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  NAND2_X1  g439(.A1(new_n354), .A2(new_n355), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n488), .B1(new_n502), .B2(new_n503), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n290), .B1(new_n477), .B2(new_n488), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n525), .B2(new_n529), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n409), .A2(new_n414), .B1(new_n455), .B2(new_n445), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n614), .A2(new_n356), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT98), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n298), .A2(new_n361), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n621), .B(KEYINPUT39), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n643), .A2(KEYINPUT40), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n643), .B2(new_n644), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n636), .B(new_n639), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G143), .ZN(G45));
  NOR2_X1   g462(.A1(new_n581), .A2(new_n622), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n620), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  NAND2_X1  g465(.A1(new_n281), .A2(new_n282), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n652), .A2(new_n277), .B1(new_n295), .B2(new_n247), .ZN(new_n653));
  OAI21_X1  g467(.A(G469), .B1(new_n653), .B2(G902), .ZN(new_n654));
  INV_X1    g468(.A(new_n360), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n655), .A3(new_n293), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n591), .A2(new_n530), .A3(new_n563), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT41), .B(G113), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G15));
  NAND4_X1  g474(.A1(new_n530), .A2(new_n604), .A3(new_n656), .A4(new_n563), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NAND4_X1  g476(.A1(new_n530), .A2(new_n656), .A3(new_n463), .A4(new_n619), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  AND4_X1   g478(.A1(new_n655), .A2(new_n654), .A3(new_n293), .A4(new_n461), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n637), .B(new_n356), .C1(new_n572), .C2(new_n573), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT101), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n584), .A2(new_n668), .A3(new_n637), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n528), .B2(new_n290), .ZN(new_n672));
  INV_X1    g486(.A(new_n512), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n522), .A2(new_n519), .B1(new_n482), .B2(new_n489), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n527), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n672), .A2(new_n562), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n665), .A2(new_n670), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G122), .ZN(G24));
  NOR3_X1   g492(.A1(new_n614), .A2(new_n672), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n649), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n656), .A2(new_n584), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n329), .ZN(G27));
  AOI21_X1  g497(.A(new_n583), .B1(new_n354), .B2(new_n355), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n530), .A2(new_n563), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(G469), .B1(new_n296), .B2(G902), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n360), .B(new_n581), .C1(new_n686), .C2(new_n293), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n621), .A4(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n687), .A2(new_n530), .A3(new_n563), .A4(new_n684), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(new_n622), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n196), .ZN(G33));
  AOI21_X1  g507(.A(new_n360), .B1(new_n686), .B2(new_n293), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n685), .A2(new_n623), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n188), .ZN(G36));
  INV_X1    g510(.A(new_n684), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n609), .A2(new_n618), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n587), .A2(new_n588), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(KEYINPUT43), .A3(new_n415), .ZN(new_n702));
  INV_X1    g516(.A(new_n415), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n415), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n704), .A2(new_n700), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n702), .B1(KEYINPUT43), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n697), .B1(new_n709), .B2(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n699), .A2(new_n708), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n278), .A2(new_n283), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n296), .A2(KEYINPUT45), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(G469), .ZN(new_n718));
  NAND2_X1  g532(.A1(G469), .A2(G902), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(KEYINPUT46), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n293), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(KEYINPUT102), .A3(new_n293), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n718), .A2(new_n719), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n723), .B(new_n724), .C1(KEYINPUT46), .C2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n726), .A2(new_n655), .A3(new_n641), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n710), .A2(new_n713), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G137), .ZN(G39));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n655), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n655), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n530), .A2(new_n563), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n649), .A3(new_n684), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G140), .ZN(G42));
  AND3_X1   g551(.A1(new_n599), .A2(new_n455), .A3(new_n445), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n530), .A2(new_n298), .A3(new_n361), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n672), .A2(new_n675), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n687), .A2(new_n740), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n614), .B(new_n697), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n695), .B1(new_n742), .B2(new_n621), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n357), .A2(new_n461), .A3(new_n589), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n569), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n565), .B2(new_n746), .ZN(new_n747));
  OAI221_X1 g561(.A(KEYINPUT106), .B1(new_n464), .B2(new_n564), .C1(new_n569), .C2(new_n745), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n657), .A2(new_n661), .A3(new_n677), .A4(new_n663), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n688), .B2(new_n691), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n703), .A2(new_n456), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n357), .A2(new_n461), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n357), .A2(new_n756), .A3(new_n461), .A4(new_n753), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n570), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n615), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n743), .A2(new_n749), .A3(new_n751), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n615), .A2(new_n758), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n747), .B2(new_n748), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT108), .A3(new_n751), .A4(new_n743), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n620), .B1(new_n623), .B2(new_n649), .ZN(new_n767));
  INV_X1    g581(.A(new_n682), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n618), .A2(new_n622), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n670), .A2(new_n634), .A3(new_n694), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n766), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n771), .B(KEYINPUT109), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(KEYINPUT52), .A3(new_n768), .A4(new_n767), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n762), .A2(new_n765), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n743), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n751), .A2(KEYINPUT112), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n776), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n774), .A2(new_n786), .A3(new_n776), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n751), .B2(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n785), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n781), .A2(new_n782), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n762), .A2(new_n765), .A3(new_n787), .A4(new_n788), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n789), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n762), .A2(new_n765), .A3(new_n777), .A4(new_n779), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT54), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n781), .A2(new_n791), .A3(KEYINPUT113), .A4(new_n782), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n794), .A2(new_n799), .A3(new_n803), .A4(new_n800), .ZN(new_n804));
  INV_X1    g618(.A(new_n656), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n697), .ZN(new_n806));
  INV_X1    g620(.A(new_n458), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n563), .A2(new_n806), .A3(new_n807), .A4(new_n635), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n808), .A2(new_n703), .A3(new_n701), .ZN(new_n809));
  INV_X1    g623(.A(new_n676), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n708), .A2(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n708), .A2(new_n813), .A3(new_n807), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n628), .A2(new_n805), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n583), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n583), .A4(new_n816), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n809), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n812), .A2(new_n814), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n806), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n679), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n654), .A2(new_n293), .ZN(new_n825));
  INV_X1    g639(.A(new_n361), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n732), .A2(new_n733), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n676), .A3(new_n684), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n821), .B(new_n824), .C1(new_n829), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n815), .A2(new_n584), .A3(new_n656), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n830), .B(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n828), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT51), .A3(new_n824), .A4(new_n821), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n822), .A2(new_n806), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n564), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n808), .A2(new_n589), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(G952), .A3(new_n274), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n564), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n823), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n840), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n841), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n840), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n835), .A2(new_n836), .A3(new_n839), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n802), .A2(new_n804), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n802), .A2(new_n854), .A3(new_n857), .A4(new_n804), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT120), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n707), .A2(new_n562), .A3(new_n583), .A4(new_n826), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT105), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n825), .B(KEYINPUT49), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n635), .A3(new_n629), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n865), .ZN(G75));
  AND2_X1   g680(.A1(new_n781), .A2(new_n791), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n290), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT56), .B1(new_n868), .B2(G210), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n327), .B(new_n337), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  NOR2_X1   g685(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n869), .B(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n274), .A2(G952), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(G51));
  XNOR2_X1  g690(.A(new_n867), .B(new_n782), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n719), .B(KEYINPUT57), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n289), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n867), .A2(new_n290), .A3(new_n718), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(G54));
  NAND3_X1  g696(.A1(new_n868), .A2(KEYINPUT58), .A3(G475), .ZN(new_n883));
  INV_X1    g697(.A(new_n403), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n883), .A2(KEYINPUT122), .A3(new_n884), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n875), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(G60));
  INV_X1    g704(.A(new_n875), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n585), .A2(new_n586), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(G478), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT59), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n877), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n802), .B2(new_n804), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n891), .B(new_n897), .C1(new_n898), .C2(new_n893), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(G63));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n867), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n891), .B1(new_n903), .B2(new_n549), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n612), .B2(new_n903), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g720(.A(new_n274), .B1(new_n332), .B2(new_n459), .ZN(new_n907));
  INV_X1    g721(.A(new_n764), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(new_n750), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n274), .ZN(new_n910));
  INV_X1    g724(.A(G898), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n327), .B1(new_n911), .B2(G953), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n910), .B(new_n912), .ZN(G69));
  INV_X1    g727(.A(new_n769), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n727), .A2(new_n846), .A3(new_n670), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n736), .A2(new_n728), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n692), .A2(new_n695), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n274), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n274), .A2(G900), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n395), .A2(new_n397), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n517), .B(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(KEYINPUT124), .A3(new_n919), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n736), .A2(new_n728), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n752), .A2(new_n581), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n643), .A2(new_n644), .A3(new_n685), .A4(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n647), .A2(KEYINPUT62), .A3(new_n914), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT62), .B1(new_n647), .B2(new_n914), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n931), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n274), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT123), .B1(new_n937), .B2(new_n924), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n939), .B(new_n925), .C1(new_n936), .C2(new_n274), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT125), .B1(new_n930), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n927), .A2(new_n929), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n937), .A2(new_n924), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n927), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT126), .B1(new_n948), .B2(new_n928), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n950), .B(new_n929), .C1(new_n927), .C2(new_n947), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n943), .A2(new_n946), .B1(new_n949), .B2(new_n951), .ZN(G72));
  NAND2_X1  g766(.A1(new_n518), .A2(new_n476), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n916), .A2(new_n909), .A3(new_n917), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI211_X1 g770(.A(new_n953), .B(new_n488), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n936), .B2(new_n909), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n875), .B(new_n957), .C1(new_n631), .C2(new_n958), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n504), .B(KEYINPUT127), .Z(new_n960));
  OAI211_X1 g774(.A(new_n798), .B(new_n956), .C1(new_n522), .C2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(G57));
endmodule


