//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(G141gat), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT78), .B1(new_n210), .B2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT79), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n211), .A2(new_n218), .A3(G141gat), .A4(new_n212), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n216), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G141gat), .B(G148gat), .Z(new_n223));
  AOI211_X1 g022(.A(new_n204), .B(new_n206), .C1(new_n223), .C2(new_n205), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  INV_X1    g026(.A(G120gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT1), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G113gat), .A2(G120gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G113gat), .B2(G120gat), .ZN(new_n233));
  AND2_X1   g032(.A1(G113gat), .A2(G120gat), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n234), .A3(G127gat), .ZN(new_n235));
  OAI21_X1  g034(.A(G134gat), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT69), .B(G127gat), .C1(new_n233), .C2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(G127gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n229), .A2(new_n238), .A3(new_n230), .ZN(new_n239));
  INV_X1    g038(.A(G134gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n222), .A2(new_n225), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n236), .A2(KEYINPUT80), .A3(new_n241), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n214), .B1(new_n250), .B2(G141gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n219), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT79), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n224), .B1(new_n255), .B2(new_n208), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n247), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n207), .B1(new_n253), .B2(new_n254), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(new_n263), .B2(new_n224), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n222), .A2(new_n265), .A3(new_n225), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n237), .A2(new_n240), .A3(new_n239), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n240), .B1(new_n237), .B2(new_n239), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n267), .A2(new_n268), .A3(new_n244), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT80), .B1(new_n236), .B2(new_n241), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n243), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n256), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n258), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT81), .A2(KEYINPUT5), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT4), .B1(new_n256), .B2(new_n242), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n267), .A2(new_n268), .ZN(new_n281));
  NOR4_X1   g080(.A1(new_n263), .A2(new_n281), .A3(new_n273), .A4(new_n224), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(new_n258), .A3(new_n272), .A4(new_n277), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n262), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G1gat), .B(G29gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT0), .ZN(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n285), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n285), .B2(new_n289), .ZN(new_n293));
  INV_X1    g092(.A(new_n289), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n294), .B(new_n262), .C1(new_n279), .C2(new_n284), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  INV_X1    g097(.A(G169gat), .ZN(new_n299));
  INV_X1    g098(.A(G176gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT65), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n304));
  AND2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n300), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT66), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n312), .A2(new_n314), .A3(new_n317), .A4(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n309), .B1(new_n310), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n318), .B2(new_n319), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n324), .A2(KEYINPUT67), .A3(new_n314), .A4(new_n312), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n298), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G183gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n329), .A3(new_n319), .ZN(new_n330));
  NOR2_X1   g129(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n333), .A2(new_n327), .A3(new_n329), .A4(new_n319), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n305), .B1(new_n306), .B2(KEYINPUT26), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n301), .A2(new_n303), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT26), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n315), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n323), .A2(KEYINPUT64), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n323), .A2(KEYINPUT64), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n311), .A3(new_n320), .A4(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT25), .B1(new_n343), .B2(KEYINPUT23), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n308), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n297), .B1(new_n326), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n304), .A2(new_n308), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n321), .A2(new_n310), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n325), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT25), .ZN(new_n353));
  INV_X1    g152(.A(new_n315), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n332), .B2(new_n334), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n355), .A2(new_n338), .B1(new_n342), .B2(new_n345), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT75), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT22), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT73), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(new_n361), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  XNOR2_X1  g166(.A(G197gat), .B(G204gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G211gat), .B(G218gat), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n372), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n373), .A3(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n353), .A2(new_n356), .ZN(new_n380));
  INV_X1    g179(.A(new_n359), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT76), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n383), .B(new_n359), .C1(new_n353), .C2(new_n356), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n349), .A3(new_n359), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT75), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT75), .B1(new_n353), .B2(new_n356), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n378), .B(new_n387), .C1(new_n390), .C2(new_n359), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n400), .A3(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G228gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n371), .B2(new_n373), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n265), .B1(new_n407), .B2(KEYINPUT83), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(KEYINPUT83), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n256), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n378), .B1(new_n349), .B2(new_n266), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n263), .B2(new_n224), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n264), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n266), .A2(new_n349), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n379), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n222), .A2(new_n225), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n407), .A2(KEYINPUT83), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(new_n408), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n405), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n412), .A2(new_n415), .ZN(new_n426));
  OAI21_X1  g225(.A(G22gat), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  NAND4_X1  g230(.A1(new_n421), .A2(new_n427), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n421), .A2(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n424), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n434), .A2(new_n406), .B1(new_n418), .B2(new_n416), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n428), .B1(new_n435), .B2(new_n420), .ZN(new_n436));
  INV_X1    g235(.A(new_n431), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n296), .A2(new_n402), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT36), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n242), .B1(new_n326), .B2(new_n347), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n353), .A2(new_n356), .A3(new_n281), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G227gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n404), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT34), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n447), .A2(KEYINPUT72), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n447), .B2(KEYINPUT72), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT70), .ZN(new_n453));
  XNOR2_X1  g252(.A(G71gat), .B(G99gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n445), .A3(new_n442), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT32), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT33), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT71), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n455), .B2(KEYINPUT33), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n451), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n459), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT71), .B1(new_n465), .B2(new_n455), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n467), .B(new_n456), .C1(new_n457), .C2(new_n459), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n447), .A2(KEYINPUT72), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT34), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n447), .A2(KEYINPUT72), .A3(new_n448), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n440), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n451), .A3(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(KEYINPUT36), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n439), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT39), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n259), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n289), .B(KEYINPUT85), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n257), .B2(new_n259), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n259), .B2(new_n482), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n481), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(KEYINPUT86), .B(new_n481), .C1(new_n487), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n487), .A2(new_n489), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(KEYINPUT40), .B1(new_n285), .B2(new_n485), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n494), .A2(new_n401), .A3(new_n399), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n392), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n386), .A2(KEYINPUT37), .A3(new_n391), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n397), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT38), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n397), .B1(new_n386), .B2(new_n391), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n395), .B1(new_n392), .B2(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n360), .A2(new_n385), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n378), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n387), .B1(new_n390), .B2(new_n359), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n498), .B1(new_n507), .B2(new_n379), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT38), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n503), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n279), .A2(new_n284), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n261), .A3(new_n485), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(new_n290), .C1(new_n289), .C2(new_n285), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n502), .A2(new_n510), .A3(new_n292), .A4(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n438), .A2(new_n432), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n480), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n296), .A2(new_n402), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n438), .B(new_n432), .C1(new_n464), .C2(new_n474), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT35), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT35), .B1(new_n513), .B2(new_n292), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n476), .A2(new_n477), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n521), .A2(new_n515), .A3(new_n402), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  INV_X1    g330(.A(G15gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(G22gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n420), .A2(G15gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT89), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n420), .A2(G15gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT16), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  INV_X1    g342(.A(new_n539), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n538), .B1(new_n536), .B2(new_n537), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n543), .B(G1gat), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(G1gat), .B1(new_n540), .B2(new_n543), .ZN(new_n548));
  OAI21_X1  g347(.A(G8gat), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(new_n543), .ZN(new_n550));
  INV_X1    g349(.A(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G8gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n546), .A4(new_n542), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G29gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n559));
  INV_X1    g358(.A(G36gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n558), .B2(KEYINPUT14), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT14), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(G29gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n559), .C1(new_n561), .C2(new_n563), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(KEYINPUT17), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n570), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT88), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n554), .A3(KEYINPUT91), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n557), .A2(new_n571), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n555), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n567), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT88), .B1(new_n567), .B2(new_n570), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n549), .A2(new_n554), .A3(KEYINPUT92), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n579), .A2(new_n587), .A3(KEYINPUT93), .A4(new_n580), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n580), .B(KEYINPUT13), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n582), .A2(new_n586), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n574), .A2(new_n576), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n595), .B1(new_n598), .B2(new_n587), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n579), .A2(new_n587), .A3(KEYINPUT18), .A4(new_n580), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n531), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(KEYINPUT94), .ZN(new_n606));
  INV_X1    g405(.A(new_n531), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n593), .A3(new_n600), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT97), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT7), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n585), .A2(new_n621), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n577), .A2(new_n571), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n623), .A2(new_n625), .A3(new_n319), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n319), .B1(new_n623), .B2(new_n625), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n363), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n577), .A2(new_n571), .A3(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n597), .B2(new_n624), .ZN(new_n631));
  OAI21_X1  g430(.A(G190gat), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n625), .A3(new_n319), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n632), .A2(G218gat), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n634), .A3(KEYINPUT96), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n628), .A2(new_n634), .A3(KEYINPUT96), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G134gat), .B(G162gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(new_n641), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G57gat), .ZN(new_n646));
  INV_X1    g445(.A(G64gat), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT95), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n646), .B2(KEYINPUT95), .ZN(new_n649));
  INV_X1    g448(.A(G71gat), .ZN(new_n650));
  INV_X1    g449(.A(G78gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT9), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n648), .B(new_n649), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n646), .A2(new_n647), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT21), .ZN(new_n661));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G127gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(KEYINPUT21), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n596), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n202), .ZN(new_n669));
  XOR2_X1   g468(.A(G183gat), .B(G211gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n667), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n613), .B2(new_n617), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n654), .B(new_n659), .C1(new_n611), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT97), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n610), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT99), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n660), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n619), .B2(new_n620), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n679), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n611), .A2(new_n677), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n687), .A2(new_n660), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n683), .A2(new_n685), .A3(new_n686), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n660), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n675), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n683), .A2(new_n685), .A3(new_n690), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(G230gat), .A3(G233gat), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(G120gat), .B(G148gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(G176gat), .B(G204gat), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n698), .B(new_n699), .Z(new_n700));
  OR2_X1    g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n691), .A2(new_n692), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n674), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n696), .A2(KEYINPUT100), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n696), .B2(KEYINPUT100), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n645), .A2(new_n673), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n525), .A2(new_n609), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n296), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT102), .B(G1gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1324gat));
  INV_X1    g514(.A(new_n402), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT16), .B(G8gat), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT103), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(G8gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(G1325gat));
  NAND3_X1  g522(.A1(new_n711), .A2(new_n532), .A3(new_n522), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n711), .A2(new_n479), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n532), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT104), .Z(G1326gat));
  INV_X1    g526(.A(new_n515), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT43), .B(G22gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1327gat));
  AOI22_X1  g530(.A1(new_n480), .A2(new_n516), .B1(new_n520), .B2(new_n523), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n637), .A2(new_n641), .A3(new_n639), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n641), .B1(new_n637), .B2(new_n639), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n609), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n672), .A3(new_n709), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(G29gat), .A3(new_n296), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT45), .Z(new_n741));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n525), .B2(new_n645), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n743), .B(new_n735), .C1(new_n517), .C2(new_n524), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n738), .B(KEYINPUT105), .Z(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n712), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n741), .B1(new_n558), .B2(new_n748), .ZN(G1328gat));
  NOR3_X1   g548(.A1(new_n739), .A2(G36gat), .A3(new_n402), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n716), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G36gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(G1329gat));
  INV_X1    g555(.A(new_n522), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n739), .A2(G43gat), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n745), .A2(new_n479), .A3(new_n746), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(G43gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g560(.A(new_n743), .B1(new_n732), .B2(new_n735), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n525), .A2(KEYINPUT44), .A3(new_n645), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n728), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  OR3_X1    g565(.A1(new_n739), .A2(G50gat), .A3(new_n515), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT107), .B1(new_n764), .B2(G50gat), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(KEYINPUT48), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n767), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n770), .A2(KEYINPUT48), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(new_n776), .ZN(G1331gat));
  NAND2_X1  g576(.A1(new_n737), .A2(new_n709), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n778), .A2(new_n673), .A3(new_n645), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n525), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n296), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT110), .B(G57gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(KEYINPUT111), .A3(new_n525), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n786), .A2(new_n716), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  NAND4_X1  g591(.A1(new_n786), .A2(G71gat), .A3(new_n479), .A4(new_n787), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n650), .B1(new_n781), .B2(new_n757), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT50), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1334gat));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n728), .A3(new_n787), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT112), .B(G78gat), .Z(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(G1335gat));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT113), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n672), .B1(KEYINPUT113), .B2(new_n801), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n737), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n736), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n736), .B2(new_n805), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n712), .A3(new_n709), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n778), .A2(new_n672), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n745), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n712), .A2(G85gat), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n810), .A2(new_n615), .B1(new_n812), .B2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n763), .A2(new_n762), .A3(new_n716), .A4(new_n811), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n616), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n745), .A2(KEYINPUT115), .A3(new_n716), .A4(new_n811), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n709), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(new_n402), .A3(G92gat), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n809), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n808), .ZN(new_n825));
  XOR2_X1   g624(.A(new_n822), .B(KEYINPUT114), .Z(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n806), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n816), .A2(G92gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n818), .A2(new_n819), .B1(new_n809), .B2(new_n822), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(new_n829), .C1(new_n833), .C2(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1337gat));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n522), .A3(new_n709), .ZN(new_n836));
  INV_X1    g635(.A(G99gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n475), .B2(new_n478), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n836), .A2(new_n837), .B1(new_n812), .B2(new_n838), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n745), .A2(new_n728), .A3(new_n811), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT117), .B(G106gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n840), .A2(new_n841), .B1(new_n842), .B2(KEYINPUT53), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n515), .A2(G106gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n809), .A2(new_n709), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n842), .A2(KEYINPUT53), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(G1339gat));
  NAND4_X1  g647(.A1(new_n735), .A2(new_n737), .A3(new_n672), .A4(new_n821), .ZN(new_n849));
  INV_X1    g648(.A(new_n675), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n703), .B(KEYINPUT54), .C1(new_n850), .C2(new_n702), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n700), .B1(new_n693), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n707), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n853), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n605), .B2(new_n608), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n598), .A2(new_n587), .A3(new_n595), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n580), .B1(new_n579), .B2(new_n587), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n530), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n608), .A2(new_n709), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n645), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n608), .A2(new_n862), .A3(new_n857), .A4(new_n855), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n733), .B2(new_n734), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n673), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n849), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n296), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n519), .A2(new_n716), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n609), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n737), .A2(new_n227), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n872), .B2(new_n709), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n821), .A2(new_n228), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  NOR2_X1   g682(.A1(new_n875), .A2(new_n673), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT120), .ZN(new_n885));
  AOI21_X1  g684(.A(G127gat), .B1(new_n884), .B2(KEYINPUT120), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n673), .A2(new_n238), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n885), .A2(new_n886), .B1(new_n878), .B2(new_n887), .ZN(G1342gat));
  XOR2_X1   g687(.A(KEYINPUT69), .B(G134gat), .Z(new_n889));
  NAND4_X1  g688(.A1(new_n870), .A2(new_n871), .A3(new_n645), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT56), .Z(new_n891));
  AOI21_X1  g690(.A(new_n735), .B1(new_n874), .B2(new_n877), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n240), .B2(new_n892), .ZN(G1343gat));
  INV_X1    g692(.A(G141gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n712), .A2(new_n402), .A3(new_n478), .A4(new_n475), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n868), .A2(KEYINPUT57), .A3(new_n728), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT57), .B1(new_n868), .B2(new_n728), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n868), .A2(new_n899), .A3(KEYINPUT57), .A4(new_n728), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n895), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(new_n609), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n479), .A2(new_n515), .A3(new_n716), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n870), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G141gat), .A3(new_n737), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT58), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n905), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n737), .B(new_n895), .C1(new_n898), .C2(new_n900), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n894), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n709), .A2(new_n250), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n904), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n250), .C1(new_n901), .C2(new_n709), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n895), .B(KEYINPUT123), .Z(new_n918));
  INV_X1    g717(.A(new_n896), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n709), .B(new_n918), .C1(new_n919), .C2(new_n897), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n915), .B1(new_n916), .B2(new_n921), .ZN(G1345gat));
  INV_X1    g721(.A(new_n904), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n202), .A3(new_n672), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n901), .A2(new_n672), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n202), .ZN(G1346gat));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n203), .A3(new_n645), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n901), .A2(new_n645), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n203), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n869), .A2(new_n712), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n519), .A2(new_n402), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n737), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(new_n299), .ZN(G1348gat));
  NOR2_X1   g733(.A1(new_n932), .A2(new_n821), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(new_n300), .ZN(G1349gat));
  AND2_X1   g735(.A1(new_n327), .A2(new_n329), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n932), .A2(new_n937), .A3(new_n673), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n318), .B1(new_n932), .B2(new_n673), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1350gat));
  NOR2_X1   g742(.A1(new_n932), .A2(new_n735), .ZN(new_n944));
  NAND2_X1  g743(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g745(.A(KEYINPUT61), .B(G190gat), .Z(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n944), .B2(new_n947), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n479), .A2(new_n712), .A3(new_n402), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n897), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n737), .B(new_n950), .C1(new_n951), .C2(new_n896), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n479), .A2(new_n515), .A3(new_n402), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  NAND2_X1  g755(.A1(new_n930), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n609), .A2(new_n953), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT125), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  OAI221_X1 g760(.A(new_n961), .B1(new_n957), .B2(new_n958), .C1(new_n952), .C2(new_n953), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n821), .A2(G204gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n930), .A2(new_n956), .A3(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n930), .A2(KEYINPUT126), .A3(new_n956), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n964), .B1(new_n970), .B2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n968), .A2(KEYINPUT127), .A3(new_n973), .A4(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n709), .B1(new_n919), .B2(new_n897), .ZN(new_n975));
  OAI21_X1  g774(.A(G204gat), .B1(new_n975), .B2(new_n950), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(G1353gat));
  INV_X1    g776(.A(new_n957), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(new_n362), .A3(new_n672), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n950), .B1(new_n951), .B2(new_n896), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n672), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n981), .B2(G211gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n363), .A3(new_n645), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n980), .A2(new_n645), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n363), .ZN(G1355gat));
endmodule


