//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n620, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n462));
  AOI211_X1 g037(.A(new_n461), .B(new_n462), .C1(new_n454), .C2(G2106), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(KEYINPUT67), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n483), .A2(new_n464), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n475), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n487), .A2(G124), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND4_X1  g068(.A1(new_n476), .A2(new_n478), .A3(G138), .A4(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(G138), .A3(new_n464), .A4(new_n496), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(new_n464), .B2(G114), .ZN(new_n502));
  NOR2_X1   g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT69), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n475), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  INV_X1    g082(.A(new_n503), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n476), .A2(new_n478), .A3(G126), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n504), .A2(new_n509), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n500), .A2(new_n501), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n507), .B1(new_n506), .B2(new_n508), .ZN(new_n514));
  NOR3_X1   g089(.A1(new_n502), .A2(KEYINPUT69), .A3(new_n503), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n498), .A2(new_n499), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(G164));
  NAND2_X1  g094(.A1(KEYINPUT73), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n524), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(G50), .A2(new_n535), .B1(new_n537), .B2(G88), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n529), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND3_X1  g115(.A1(new_n533), .A2(G51), .A3(G543), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n533), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n544));
  INV_X1    g119(.A(new_n524), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  XOR2_X1   g122(.A(KEYINPUT77), .B(G90), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n537), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT76), .B(G52), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n535), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n552), .B1(new_n549), .B2(new_n551), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  XNOR2_X1  g135(.A(KEYINPUT79), .B(G81), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n533), .A2(new_n524), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G43), .ZN(new_n564));
  OAI221_X1 g139(.A(new_n562), .B1(new_n563), .B2(new_n526), .C1(new_n534), .C2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G860), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n545), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n537), .A2(G91), .B1(new_n575), .B2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n535), .A2(KEYINPUT9), .A3(G53), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n534), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(G299));
  OR2_X1    g156(.A1(new_n524), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n537), .A2(G87), .B1(G651), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n534), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n535), .A2(KEYINPUT80), .A3(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n545), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n535), .A2(G48), .B1(new_n591), .B2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n537), .A2(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n537), .A2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n535), .A2(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n595), .B(new_n596), .C1(new_n526), .C2(new_n597), .ZN(G290));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n536), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT10), .B1(new_n536), .B2(new_n599), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n545), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n535), .A2(G54), .B1(new_n605), .B2(G651), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n602), .A2(KEYINPUT81), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n600), .A3(new_n601), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G284));
  OAI21_X1  g189(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  NAND2_X1  g190(.A1(G299), .A2(new_n612), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n565), .B(new_n622), .S(G868), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n487), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G135), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n674), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT83), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(G229));
  MUX2_X1   g259(.A(G24), .B(G290), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT84), .Z(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n487), .A2(G119), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n484), .A2(G131), .ZN(new_n691));
  OR2_X1    g266(.A1(G95), .A2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NOR4_X1   g273(.A1(new_n688), .A2(new_n689), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT85), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n700), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1971), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n703), .B(KEYINPUT85), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(new_n705), .ZN(new_n712));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n707), .A2(new_n710), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n699), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT36), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n722), .B(new_n699), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G299), .A2(G16), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n700), .A2(KEYINPUT23), .A3(G20), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n727));
  INV_X1    g302(.A(G20), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G16), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G1956), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n700), .A2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G168), .B2(new_n700), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT86), .B1(G4), .B2(G16), .ZN(new_n745));
  OR3_X1    g320(.A1(KEYINPUT86), .A2(G4), .A3(G16), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n745), .B(new_n746), .C1(new_n611), .C2(new_n700), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1348), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n487), .A2(G129), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n484), .A2(G141), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  NAND4_X1  g329(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G32), .B(new_n757), .S(G29), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT27), .B(G1996), .Z(new_n759));
  NOR3_X1   g334(.A1(new_n758), .A2(KEYINPUT91), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n743), .B2(new_n742), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n749), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n763));
  INV_X1    g338(.A(G26), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n484), .A2(G140), .ZN(new_n768));
  NOR2_X1   g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT88), .Z(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n766), .B1(new_n772), .B2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n765), .B1(new_n773), .B2(new_n763), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT94), .B(G28), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT30), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n780), .C1(new_n629), .C2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT95), .ZN(new_n782));
  NOR2_X1   g357(.A1(G27), .A2(G29), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G164), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(KEYINPUT24), .A2(G34), .ZN(new_n788));
  NAND2_X1  g363(.A1(KEYINPUT24), .A2(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G160), .B2(G29), .ZN(new_n791));
  MUX2_X1   g366(.A(new_n790), .B(new_n791), .S(KEYINPUT89), .Z(new_n792));
  AOI211_X1 g367(.A(new_n775), .B(new_n787), .C1(G2084), .C2(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(G2084), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n758), .A2(new_n759), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n700), .A2(G19), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n565), .B2(G16), .ZN(new_n797));
  MUX2_X1   g372(.A(new_n796), .B(new_n797), .S(KEYINPUT87), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1341), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G2072), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT25), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(new_n464), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n803), .B(new_n805), .C1(new_n484), .C2(G139), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G29), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G29), .B2(G33), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n740), .A2(new_n741), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT91), .B1(new_n758), .B2(new_n759), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n793), .A2(new_n800), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n774), .A2(G2067), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n801), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n762), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n724), .A2(new_n732), .A3(new_n737), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n779), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n779), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT29), .B(G2090), .Z(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  NOR2_X1   g395(.A1(new_n816), .A2(new_n820), .ZN(G311));
  NOR3_X1   g396(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n822), .A2(new_n761), .A3(new_n749), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n721), .B2(new_n723), .ZN(new_n824));
  INV_X1    g399(.A(new_n820), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n824), .A2(new_n825), .A3(new_n732), .A4(new_n737), .ZN(G150));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(G55), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n533), .A2(G543), .A3(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n828), .B1(new_n829), .B2(new_n526), .C1(new_n536), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n565), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n831), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n535), .A2(G43), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n563), .A2(new_n526), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT98), .A4(new_n562), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n565), .A2(new_n831), .A3(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n619), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n566), .B1(new_n845), .B2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n833), .B1(new_n848), .B2(new_n849), .ZN(G145));
  NAND2_X1  g425(.A1(new_n500), .A2(new_n511), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n772), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n484), .A2(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n464), .A2(G118), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT100), .Z(new_n856));
  OAI21_X1  g431(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G130), .B2(new_n487), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n632), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G160), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n492), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n492), .A2(new_n862), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n629), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(G162), .A2(G160), .ZN(new_n867));
  INV_X1    g442(.A(new_n629), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n863), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n694), .B(KEYINPUT101), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n866), .B2(new_n869), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n755), .A2(new_n806), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n757), .B2(new_n806), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n866), .A2(new_n869), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n870), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n880), .B2(new_n872), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n861), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n878), .A3(new_n872), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n860), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n622), .B(new_n842), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n608), .A2(new_n576), .A3(new_n580), .A4(new_n577), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n602), .A2(G299), .A3(new_n606), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n892), .B2(new_n891), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(KEYINPUT103), .A3(new_n895), .ZN(new_n899));
  XNOR2_X1  g474(.A(G299), .B(new_n608), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n894), .B2(KEYINPUT41), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n898), .B(new_n899), .C1(new_n889), .C2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n702), .B(KEYINPUT104), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(G290), .B(G305), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G303), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(G303), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n904), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n903), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n903), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n836), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n836), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  INV_X1    g496(.A(new_n900), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  AND3_X1   g499(.A1(G286), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(G286), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n842), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G168), .A2(KEYINPUT105), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(new_n558), .C1(new_n553), .C2(new_n554), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n840), .B(new_n841), .C1(new_n926), .C2(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n928), .B2(new_n932), .ZN(new_n935));
  OAI211_X1 g510(.A(KEYINPUT41), .B(new_n922), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n930), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n913), .B(new_n936), .C1(new_n895), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n941), .B2(KEYINPUT108), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n902), .B1(new_n934), .B2(new_n935), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n894), .A3(new_n933), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n913), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT41), .B1(new_n934), .B2(new_n935), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n894), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n913), .A4(new_n936), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n942), .A2(new_n943), .A3(new_n948), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n944), .A2(new_n913), .A3(new_n945), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n883), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n921), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT107), .B1(new_n955), .B2(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n920), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n941), .A2(KEYINPUT108), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(new_n883), .A3(new_n948), .A4(new_n952), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n920), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n959), .A2(new_n968), .ZN(G397));
  AOI21_X1  g544(.A(G1384), .B1(new_n500), .B2(new_n511), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n468), .A2(new_n471), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n772), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n757), .B2(G1996), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(G1996), .B2(new_n755), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n694), .A2(new_n696), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n694), .A2(new_n696), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G290), .B(G1986), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  INV_X1    g560(.A(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n592), .A2(new_n986), .A3(new_n593), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n592), .B2(new_n593), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(KEYINPUT49), .A3(new_n987), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n469), .A2(new_n470), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n464), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n466), .A2(new_n467), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n994), .B(G40), .C1(new_n464), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n516), .B2(new_n517), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n990), .A2(new_n992), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1003), .B2(G288), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n702), .B2(G1976), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1002), .B(new_n1005), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT111), .B(G1971), .Z(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n512), .A2(new_n518), .A3(new_n997), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n996), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(new_n997), .C1(new_n516), .C2(new_n517), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n973), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT112), .B(G2090), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1000), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT55), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G303), .A2(G8), .ZN(new_n1030));
  MUX2_X1   g605(.A(new_n1027), .B(new_n1029), .S(new_n1030), .Z(new_n1031));
  AOI21_X1  g606(.A(new_n1008), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n973), .B(new_n1034), .C1(new_n1011), .C2(KEYINPUT50), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n1024), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1000), .B1(new_n1018), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1033), .B1(new_n1038), .B2(new_n1031), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1030), .A2(new_n1029), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1030), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1027), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT110), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1036), .B1(new_n1046), .B2(new_n1010), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT116), .B(new_n1042), .C1(new_n1047), .C2(new_n1000), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1032), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n512), .A2(new_n518), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(KEYINPUT117), .A3(KEYINPUT45), .A4(new_n997), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n971), .A2(new_n996), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n741), .B1(new_n1057), .B2(new_n1022), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT51), .B1(new_n1058), .B2(G168), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1000), .B1(new_n1058), .B2(G168), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  AOI221_X4 g637(.A(G286), .B1(new_n1057), .B2(new_n1022), .C1(new_n1056), .C2(new_n741), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT51), .B1(new_n1063), .B2(new_n1000), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1050), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT125), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1061), .A2(new_n1064), .A3(new_n1062), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(KEYINPUT62), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1046), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n1072), .B2(new_n785), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1023), .A2(new_n736), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1074), .B(new_n1075), .C1(new_n1056), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1067), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n999), .A2(new_n976), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT60), .B(new_n1081), .C1(new_n1022), .C2(G1348), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n619), .A3(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1022), .A2(G1348), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1081), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(KEYINPUT124), .A3(new_n611), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1035), .A2(new_n731), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT119), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1035), .A2(new_n1094), .A3(new_n731), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1013), .A2(new_n1015), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT120), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1013), .A2(new_n1099), .A3(new_n1015), .A4(new_n1096), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1093), .A2(new_n1095), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  XOR2_X1   g677(.A(G299), .B(KEYINPUT57), .Z(new_n1103));
  NAND4_X1  g678(.A1(new_n1101), .A2(KEYINPUT122), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT121), .B(G1996), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1013), .A2(new_n1015), .A3(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n996), .B2(new_n998), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n565), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1109), .B(KEYINPUT59), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(KEYINPUT122), .A3(new_n1103), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(KEYINPUT122), .A2(KEYINPUT123), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1102), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1091), .A2(new_n1104), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n611), .B1(new_n1086), .B2(new_n1081), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G301), .B(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1077), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1075), .B(KEYINPUT126), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1076), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1055), .A2(new_n1126), .ZN(new_n1127));
  OR4_X1    g702(.A1(new_n1123), .A2(new_n1073), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1080), .A2(new_n1122), .A3(new_n1124), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1049), .B1(new_n1079), .B2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1058), .A2(new_n1000), .A3(G286), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1032), .A2(new_n1039), .A3(new_n1048), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1133), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(new_n1032), .A3(KEYINPUT63), .A4(new_n1131), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1001), .B(KEYINPUT114), .Z(new_n1141));
  AND3_X1   g716(.A1(new_n1002), .A2(new_n1003), .A3(new_n702), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n988), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1008), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n984), .B1(new_n1130), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n981), .B(KEYINPUT127), .Z(new_n1149));
  AND2_X1   g724(.A1(new_n979), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n772), .A2(G2067), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n975), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n977), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n975), .B1(new_n1153), .B2(new_n755), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n974), .B2(G1996), .ZN(new_n1156));
  OR3_X1    g731(.A1(new_n974), .A2(new_n1155), .A3(G1996), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n982), .A2(new_n975), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT48), .Z(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1148), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g740(.A(G319), .B1(new_n647), .B2(new_n648), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n1167), .A2(G229), .ZN(new_n1168));
  AND2_X1   g742(.A1(new_n887), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g743(.A(new_n1169), .B(new_n663), .C1(new_n957), .C2(new_n958), .ZN(G225));
  INV_X1    g744(.A(G225), .ZN(G308));
endmodule


