//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(G116), .B(G119), .Z(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(new_n188), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT11), .A3(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G131), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(new_n199), .A3(new_n203), .A4(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n207), .A2(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(new_n210), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n205), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT30), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(G143), .B2(new_n206), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n216), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n207), .A2(new_n209), .A3(new_n222), .A4(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n200), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n196), .A2(G137), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n204), .A3(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n220), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n221), .B1(new_n220), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n194), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n220), .A2(new_n231), .A3(new_n191), .A4(new_n193), .ZN(new_n235));
  INV_X1    g049(.A(G237), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G210), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(G101), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT31), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT31), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n234), .A2(new_n244), .A3(new_n235), .A4(new_n241), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n241), .B(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n220), .A2(new_n231), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n194), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n249), .B2(new_n235), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n235), .A2(new_n247), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n246), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n243), .A2(new_n245), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(G472), .ZN(new_n256));
  INV_X1    g070(.A(G902), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n243), .A2(new_n258), .A3(new_n253), .A4(new_n245), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT32), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n250), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n263), .A2(new_n251), .A3(KEYINPUT29), .A4(new_n241), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n250), .A2(new_n252), .A3(new_n246), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n265), .A2(KEYINPUT29), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n234), .A2(new_n235), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(new_n241), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n257), .B(new_n264), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G472), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n260), .B2(new_n261), .ZN(new_n273));
  AND4_X1   g087(.A1(new_n256), .A2(new_n255), .A3(new_n257), .A4(new_n259), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G137), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n277), .B(new_n278), .Z(new_n279));
  INV_X1    g093(.A(G140), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  INV_X1    g095(.A(G125), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G140), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT69), .A3(KEYINPUT16), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT16), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n280), .A3(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n283), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n206), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n285), .A2(new_n290), .A3(G146), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G128), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT68), .B1(new_n296), .B2(KEYINPUT23), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n224), .A2(G119), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n224), .B(G119), .C1(KEYINPUT68), .C2(KEYINPUT23), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G110), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n298), .A2(new_n296), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT24), .B(G110), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n294), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  INV_X1    g120(.A(G110), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n307), .A3(new_n300), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n304), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n281), .A2(new_n283), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n281), .B2(new_n283), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n206), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n316), .A3(new_n309), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n311), .A2(new_n293), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n305), .A2(new_n306), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n306), .B1(new_n305), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n279), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n279), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n305), .A2(new_n318), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(KEYINPUT72), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n325), .A2(G902), .B1(KEYINPUT73), .B2(KEYINPUT25), .ZN(new_n326));
  INV_X1    g140(.A(G217), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(G234), .B2(new_n257), .ZN(new_n328));
  NOR2_X1   g142(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n321), .A2(new_n257), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n325), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(G902), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n187), .B1(new_n276), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n260), .A2(new_n261), .B1(new_n269), .B2(G472), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT67), .B1(new_n274), .B2(KEYINPUT32), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n260), .A2(new_n272), .A3(new_n261), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n335), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT74), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G469), .ZN(new_n343));
  INV_X1    g157(.A(G104), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G107), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G104), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT3), .B1(new_n344), .B2(G107), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n346), .A3(G104), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT75), .B(G101), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n216), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n224), .B1(new_n358), .B2(KEYINPUT78), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n223), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n226), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n348), .B(new_n367), .C1(new_n353), .C2(new_n354), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n227), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n205), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(KEYINPUT12), .B(new_n205), .C1(new_n365), .C2(new_n369), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  INV_X1    g189(.A(G227), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G953), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n375), .B(new_n377), .Z(new_n378));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n225), .B2(new_n226), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n368), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n364), .A2(new_n379), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n353), .A2(G101), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT77), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n353), .A2(new_n388), .A3(G101), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n215), .A2(new_n219), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n353), .A2(G101), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n392), .B(KEYINPUT4), .C1(new_n354), .C2(new_n353), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n366), .A2(KEYINPUT80), .A3(new_n368), .A4(new_n380), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n383), .A2(new_n384), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n378), .B1(new_n396), .B2(new_n205), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n374), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n384), .A2(new_n394), .ZN(new_n399));
  INV_X1    g213(.A(new_n205), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n399), .A2(new_n400), .A3(new_n383), .A4(new_n395), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n205), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n378), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n343), .B(new_n257), .C1(new_n398), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(G469), .A2(G902), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(new_n378), .C1(new_n396), .C2(new_n205), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n378), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n396), .A2(new_n205), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n374), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT82), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n406), .B1(new_n418), .B2(G469), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n390), .A2(new_n194), .A3(new_n393), .ZN(new_n424));
  INV_X1    g238(.A(G116), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n425), .A2(KEYINPUT5), .A3(G119), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n427), .A2(G113), .B1(new_n189), .B2(new_n190), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n366), .A2(new_n428), .A3(new_n368), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G122), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n424), .A2(new_n429), .A3(new_n431), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n282), .B1(new_n215), .B2(new_n219), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n225), .A2(new_n282), .A3(new_n226), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n237), .A2(G224), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n430), .A2(new_n442), .A3(new_n432), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n435), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT83), .B1(new_n428), .B2(new_n356), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n446));
  INV_X1    g260(.A(new_n426), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(G113), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n191), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n355), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n429), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n431), .B(KEYINPUT8), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n440), .A2(KEYINPUT7), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n436), .B2(new_n438), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n452), .A2(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n439), .A2(KEYINPUT7), .A3(new_n440), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n456), .A2(new_n454), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n457), .A2(new_n434), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n257), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n423), .B1(new_n444), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n435), .A2(new_n441), .A3(new_n443), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n463), .A2(new_n257), .A3(new_n422), .A4(new_n460), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n421), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G234), .A2(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G952), .A3(new_n237), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT87), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(G902), .A3(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n313), .B2(new_n314), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n289), .A2(KEYINPUT19), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n206), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT86), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n236), .A2(new_n237), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n208), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n236), .A2(new_n237), .A3(G143), .A4(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G131), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n203), .A3(new_n481), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n475), .A2(new_n486), .A3(new_n206), .A4(new_n476), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n478), .A2(new_n485), .A3(new_n293), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n480), .A2(KEYINPUT85), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n315), .B1(new_n206), .B2(new_n284), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n344), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n483), .A2(new_n499), .A3(new_n484), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n482), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n292), .A2(new_n500), .A3(new_n293), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n493), .A3(new_n496), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n505));
  INV_X1    g319(.A(G475), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n257), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n496), .B1(new_n488), .B2(new_n493), .ZN(new_n508));
  INV_X1    g322(.A(new_n503), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n506), .B(new_n257), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n496), .B1(new_n502), .B2(new_n493), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n257), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n507), .A2(new_n511), .B1(G475), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G128), .B(G143), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT13), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n208), .A2(G128), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(G134), .C1(KEYINPUT13), .C2(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(G116), .B(G122), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G107), .ZN(new_n520));
  XNOR2_X1  g334(.A(G116), .B(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n346), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n196), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n515), .B(new_n196), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n425), .A2(KEYINPUT14), .A3(G122), .ZN(new_n527));
  OAI211_X1 g341(.A(G107), .B(new_n527), .C1(new_n519), .C2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT9), .B(G234), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n531), .A2(new_n327), .A3(G953), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n529), .A3(new_n532), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n536), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n514), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n531), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NOR4_X1   g357(.A1(new_n419), .A2(new_n473), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n336), .A2(new_n342), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n354), .ZN(G3));
  NOR2_X1   g360(.A1(new_n419), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n534), .A2(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n534), .A2(KEYINPUT33), .A3(new_n535), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n550), .A2(new_n257), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n536), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n537), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT88), .B1(new_n536), .B2(G478), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n552), .A2(G478), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n507), .A2(new_n511), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n513), .A2(G475), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n473), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n260), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n547), .A2(new_n341), .A3(new_n562), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT34), .B(G104), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(G6));
  NAND2_X1  g383(.A1(new_n514), .A2(new_n539), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n473), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n547), .A2(new_n341), .A3(new_n566), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G107), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT89), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(new_n574), .ZN(G9));
  OR2_X1    g389(.A1(new_n322), .A2(KEYINPUT36), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n323), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n323), .A2(new_n576), .ZN(new_n578));
  INV_X1    g392(.A(new_n333), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT90), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n331), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n544), .A2(new_n566), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT37), .B(G110), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G12));
  NAND4_X1  g399(.A1(new_n340), .A2(new_n547), .A3(new_n465), .A4(new_n582), .ZN(new_n586));
  INV_X1    g400(.A(G900), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n469), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n468), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n570), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n224), .ZN(G30));
  XOR2_X1   g407(.A(new_n589), .B(KEYINPUT39), .Z(new_n594));
  NAND2_X1  g408(.A1(new_n547), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n595), .A2(KEYINPUT40), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n275), .A2(new_n273), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n249), .A2(new_n235), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n267), .A2(new_n241), .B1(new_n598), .B2(new_n246), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n599), .B2(G902), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n597), .A2(new_n262), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n582), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n462), .A2(new_n464), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT38), .Z(new_n604));
  NOR3_X1   g418(.A1(new_n514), .A2(new_n421), .A3(new_n540), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n595), .A2(KEYINPUT40), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n596), .A2(new_n602), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G143), .ZN(G45));
  AND3_X1   g424(.A1(new_n340), .A2(new_n547), .A3(new_n582), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT91), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n559), .ZN(new_n613));
  INV_X1    g427(.A(new_n557), .ZN(new_n614));
  INV_X1    g428(.A(new_n589), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n611), .A2(new_n612), .A3(new_n465), .A4(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT91), .B1(new_n586), .B2(new_n616), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G146), .ZN(G48));
  AND2_X1   g435(.A1(new_n396), .A2(new_n205), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n411), .B1(new_n622), .B2(new_n412), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n372), .A2(new_n373), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n401), .A3(new_n378), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n626), .A2(new_n343), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n542), .A3(new_n404), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n340), .A2(new_n341), .A3(new_n562), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT41), .B(G113), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G15));
  NAND4_X1  g446(.A1(new_n340), .A2(new_n341), .A3(new_n571), .A4(new_n629), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT92), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n335), .B1(new_n597), .B2(new_n337), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n636), .A2(KEYINPUT92), .A3(new_n571), .A4(new_n629), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G116), .ZN(G18));
  NAND2_X1  g453(.A1(new_n582), .A2(new_n465), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n628), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n541), .B1(new_n468), .B2(new_n471), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n340), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G119), .ZN(G21));
  AND3_X1   g458(.A1(new_n563), .A2(KEYINPUT95), .A3(G472), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT95), .B1(new_n563), .B2(G472), .ZN(new_n646));
  NOR2_X1   g460(.A1(G472), .A2(G902), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT93), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n243), .A2(new_n650), .A3(new_n253), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n650), .B1(new_n243), .B2(new_n253), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n649), .B1(new_n653), .B2(new_n245), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n645), .A2(new_n646), .A3(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n473), .A2(new_n540), .A3(new_n514), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n629), .A3(new_n656), .A4(new_n341), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G122), .ZN(G24));
  NAND2_X1  g472(.A1(new_n616), .A2(KEYINPUT96), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n560), .A2(new_n660), .A3(new_n615), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n641), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT97), .B(G125), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G27));
  AND3_X1   g479(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n666), .A2(KEYINPUT99), .A3(KEYINPUT32), .A4(new_n256), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n260), .B2(new_n261), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n337), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n341), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n543), .A2(new_n421), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n462), .A2(new_n464), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n410), .A2(new_n413), .A3(G469), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n405), .B(KEYINPUT98), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n626), .B2(new_n343), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n673), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n660), .B1(new_n560), .B2(new_n615), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n514), .A2(new_n557), .A3(KEYINPUT96), .A4(new_n589), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n678), .B(KEYINPUT42), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT100), .B1(new_n671), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n681), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n341), .A4(new_n670), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n340), .A2(new_n341), .A3(new_n662), .A4(new_n678), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n682), .A2(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n203), .ZN(G33));
  NAND3_X1  g503(.A1(new_n636), .A2(new_n590), .A3(new_n678), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G134), .ZN(G36));
  NAND3_X1  g505(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT45), .ZN(new_n692));
  OAI211_X1 g506(.A(G469), .B(new_n692), .C1(new_n418), .C2(KEYINPUT45), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(KEYINPUT46), .B1(new_n343), .B2(new_n626), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n695), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n675), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n543), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n565), .A2(new_n582), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT103), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n614), .A2(new_n514), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n705), .B1(KEYINPUT102), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n708));
  MUX2_X1   g522(.A(new_n705), .B(new_n707), .S(new_n708), .Z(new_n709));
  AND2_X1   g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT44), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n603), .A2(new_n421), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n710), .B2(KEYINPUT44), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n702), .A2(new_n711), .A3(new_n594), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G137), .ZN(G39));
  NAND2_X1  g530(.A1(new_n697), .A2(new_n701), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n542), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n702), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n340), .A2(new_n341), .A3(new_n713), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n617), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT104), .B(G140), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G42));
  NAND2_X1  g539(.A1(new_n627), .A2(new_n404), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n672), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n705), .B(new_n729), .C1(new_n728), .C2(new_n727), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n341), .A3(new_n604), .A4(new_n601), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n545), .A2(new_n572), .A3(new_n583), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n630), .A2(new_n643), .A3(new_n657), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n635), .B2(new_n637), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n735), .A3(new_n567), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n682), .A2(new_n685), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n686), .A2(new_n687), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n462), .A2(new_n464), .A3(new_n672), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n404), .A2(new_n674), .A3(new_n675), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n659), .B2(new_n661), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n655), .A2(new_n743), .A3(new_n744), .A4(new_n582), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n564), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n563), .A2(KEYINPUT95), .A3(G472), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n653), .A2(new_n245), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n648), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(new_n582), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT105), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n713), .A2(new_n541), .A3(new_n589), .ZN(new_n756));
  AND4_X1   g570(.A1(new_n340), .A2(new_n547), .A3(new_n582), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n739), .A2(new_n690), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n732), .B1(new_n736), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n690), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n688), .A2(new_n761), .A3(new_n754), .A4(new_n757), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n630), .A2(new_n643), .A3(new_n657), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n638), .A2(new_n567), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(KEYINPUT106), .A3(new_n733), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n663), .B1(new_n586), .B2(new_n591), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n618), .B2(new_n619), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n605), .A2(new_n603), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n589), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n602), .A2(new_n542), .A3(new_n741), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n760), .A2(new_n765), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n772), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n736), .A2(new_n759), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT54), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n760), .A3(new_n765), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  INV_X1    g601(.A(new_n468), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n709), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n655), .A2(new_n341), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n628), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n421), .A3(new_n604), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n727), .A2(new_n740), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT107), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n789), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n751), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n719), .A2(new_n721), .B1(new_n543), .B2(new_n727), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n790), .A2(new_n791), .A3(new_n713), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n795), .B(new_n801), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n797), .A2(new_n601), .A3(new_n341), .A4(new_n788), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n613), .A3(new_n614), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n702), .A2(new_n720), .ZN(new_n809));
  AOI211_X1 g623(.A(KEYINPUT47), .B(new_n543), .C1(new_n697), .C2(new_n701), .ZN(new_n810));
  OAI22_X1  g624(.A1(new_n809), .A2(new_n810), .B1(new_n542), .B2(new_n726), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n811), .A2(new_n803), .B1(new_n800), .B2(new_n799), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  INV_X1    g627(.A(new_n807), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n795), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n798), .A2(new_n671), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT48), .Z(new_n818));
  OR2_X1    g632(.A1(new_n806), .A2(new_n561), .ZN(new_n819));
  INV_X1    g633(.A(G952), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n820), .B(G953), .C1(new_n792), .C2(new_n465), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n787), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(KEYINPUT108), .B(new_n822), .C1(new_n808), .C2(new_n815), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n786), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(G952), .A2(G953), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n731), .B1(new_n826), .B2(new_n827), .ZN(G75));
  NAND2_X1  g642(.A1(new_n820), .A2(G953), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT110), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n435), .A2(new_n443), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT109), .Z(new_n832));
  XOR2_X1   g646(.A(new_n441), .B(KEYINPUT55), .Z(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n257), .B1(new_n777), .B2(new_n780), .ZN(new_n835));
  AOI211_X1 g649(.A(KEYINPUT56), .B(new_n834), .C1(new_n835), .C2(G210), .ZN(new_n836));
  INV_X1    g650(.A(new_n834), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n781), .A2(G210), .A3(G902), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n830), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT111), .B(new_n830), .C1(new_n836), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(G51));
  INV_X1    g659(.A(new_n830), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n775), .A2(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n783), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n782), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n675), .B(KEYINPUT112), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT57), .Z(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n398), .A2(new_n403), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT113), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n835), .A2(new_n694), .A3(new_n695), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n846), .B1(new_n855), .B2(new_n856), .ZN(G54));
  AND3_X1   g671(.A1(new_n835), .A2(KEYINPUT58), .A3(G475), .ZN(new_n858));
  INV_X1    g672(.A(new_n504), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n846), .B1(new_n860), .B2(new_n861), .ZN(G60));
  NAND2_X1  g676(.A1(new_n550), .A2(new_n551), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(G478), .A2(G902), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT59), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n849), .A2(KEYINPUT114), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n782), .B2(new_n785), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n846), .B1(new_n868), .B2(new_n863), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n864), .B(new_n866), .C1(new_n782), .C2(new_n848), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n867), .A2(new_n869), .A3(new_n872), .ZN(G63));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT116), .ZN(new_n877));
  XNOR2_X1  g691(.A(KEYINPUT115), .B(KEYINPUT60), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n777), .B2(new_n780), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n875), .B1(new_n881), .B2(new_n332), .ZN(new_n882));
  OAI211_X1 g696(.A(KEYINPUT118), .B(new_n325), .C1(new_n847), .C2(new_n880), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n577), .A2(new_n578), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT61), .A3(new_n830), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n874), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n889), .B(new_n846), .C1(new_n881), .C2(new_n885), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n882), .A4(new_n883), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n325), .B1(new_n847), .B2(new_n880), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n830), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n886), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n893), .B2(new_n830), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n889), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(G66));
  INV_X1    g713(.A(G224), .ZN(new_n900));
  OAI21_X1  g714(.A(G953), .B1(new_n470), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n736), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(G953), .ZN(new_n903));
  INV_X1    g717(.A(new_n832), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(G898), .B2(new_n237), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(G69));
  NOR2_X1   g720(.A1(new_n232), .A2(new_n233), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n475), .A2(new_n476), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n688), .A2(new_n761), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n723), .A2(new_n715), .A3(new_n767), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n702), .A2(new_n594), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n671), .A3(new_n769), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n915), .B2(new_n237), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n587), .B2(new_n237), .ZN(new_n917));
  OAI21_X1  g731(.A(G953), .B1(new_n376), .B2(new_n587), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n723), .A2(new_n715), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n336), .A2(new_n342), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n921), .A2(new_n595), .A3(new_n713), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n561), .A2(new_n570), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n922), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n767), .A2(new_n609), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(KEYINPUT121), .A3(KEYINPUT62), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n767), .A2(new_n936), .A3(new_n609), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT120), .Z(new_n938));
  AND3_X1   g752(.A1(new_n920), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n910), .B1(new_n939), .B2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n917), .A2(new_n919), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G72));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n920), .A2(new_n935), .A3(new_n938), .A4(new_n902), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g763(.A(new_n241), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n267), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n945), .A2(new_n952), .A3(new_n947), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n777), .A2(new_n784), .ZN(new_n955));
  INV_X1    g769(.A(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n267), .A2(new_n950), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n955), .A2(new_n956), .A3(new_n947), .A4(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n947), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n915), .B2(new_n902), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n958), .B(new_n830), .C1(new_n960), .C2(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n944), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n960), .ZN(new_n963));
  INV_X1    g777(.A(new_n957), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n846), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n949), .A2(new_n953), .A3(new_n951), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT126), .A4(new_n958), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n962), .A2(new_n967), .ZN(G57));
endmodule


