//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT22), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(G137), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT74), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n195), .A2(new_n199), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT73), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT73), .B1(new_n207), .B2(new_n208), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n202), .A2(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT75), .B(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G140), .ZN(new_n216));
  NOR2_X1   g030(.A1(G125), .A2(G140), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G140), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT75), .A2(G125), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT75), .A2(G125), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n220), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT16), .B1(new_n228), .B2(new_n217), .ZN(new_n229));
  AOI21_X1  g043(.A(G146), .B1(new_n229), .B2(new_n221), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n213), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  XOR2_X1   g046(.A(G125), .B(G140), .Z(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n201), .A2(new_n203), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n207), .A2(new_n208), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(G146), .A3(new_n221), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n231), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n232), .B1(new_n231), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n193), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n223), .B1(new_n219), .B2(new_n222), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n238), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(new_n213), .B1(new_n238), .B2(new_n237), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n193), .B1(new_n245), .B2(new_n232), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n188), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n248), .A2(new_n250), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n242), .A2(new_n247), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT77), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n189), .B(new_n251), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n241), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n232), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n246), .B1(new_n258), .B2(new_n193), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n189), .A2(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT64), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT0), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n265), .A2(new_n267), .B1(new_n268), .B2(new_n194), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n223), .A2(KEYINPUT65), .A3(G143), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT65), .B1(new_n223), .B2(G143), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n269), .A2(new_n275), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G137), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(G137), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n280), .A2(new_n283), .A3(new_n286), .A4(new_n281), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(KEYINPUT66), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n289), .A3(G131), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n288), .A2(KEYINPUT68), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT68), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n277), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n270), .B2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n223), .A2(G143), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n271), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n276), .A2(new_n301), .A3(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n281), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n279), .A2(G137), .ZN(new_n306));
  OAI21_X1  g120(.A(G131), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n287), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n293), .A2(new_n311), .A3(KEYINPUT30), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n314));
  INV_X1    g128(.A(new_n308), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n277), .A2(new_n290), .A3(new_n288), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT2), .B(G113), .Z(new_n318));
  XNOR2_X1  g132(.A(G116), .B(G119), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT31), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G210), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT27), .Z(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT26), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n320), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n293), .A2(new_n331), .A3(new_n308), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n324), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n321), .B1(new_n310), .B2(new_n312), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT31), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n320), .B1(new_n315), .B2(new_n316), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n331), .A4(new_n308), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n330), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n342), .A2(KEYINPUT70), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT70), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n335), .B(new_n337), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G472), .A2(G902), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT71), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT32), .B1(new_n346), .B2(new_n349), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n332), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n313), .B2(new_n322), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT72), .B1(new_n354), .B2(new_n330), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n343), .C1(new_n336), .C2(new_n353), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n342), .A2(new_n343), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n293), .A2(new_n308), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n320), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n339), .A2(new_n341), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n363), .A2(new_n364), .A3(new_n343), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G472), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n262), .B1(new_n352), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G104), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G107), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n329), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n370), .A3(G104), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n376), .A2(new_n373), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n372), .B2(G107), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n329), .A4(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(new_n376), .A3(new_n329), .A4(new_n373), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n374), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(new_n304), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n294), .A2(KEYINPUT81), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n298), .A2(new_n388), .A3(KEYINPUT1), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(G128), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n276), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n303), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n383), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n386), .B1(new_n383), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n288), .A2(new_n290), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n291), .A2(new_n292), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT12), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n399), .A2(KEYINPUT12), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n190), .A2(G227), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n379), .A2(new_n376), .A3(new_n373), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G101), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n381), .B(new_n378), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n277), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n383), .A2(KEYINPUT10), .A3(new_n304), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n374), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n381), .A2(KEYINPUT80), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n390), .A2(new_n391), .B1(new_n300), .B2(new_n302), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n383), .A2(new_n393), .A3(new_n386), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n414), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT84), .B1(new_n424), .B2(new_n400), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n394), .B2(new_n395), .ZN(new_n426));
  INV_X1    g240(.A(new_n414), .ZN(new_n427));
  AND4_X1   g241(.A1(KEYINPUT84), .A2(new_n426), .A3(new_n427), .A4(new_n400), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n402), .B(new_n406), .C1(new_n425), .C2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n424), .A2(new_n400), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n427), .A3(new_n400), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n424), .A2(KEYINPUT84), .A3(new_n400), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n435), .B2(new_n406), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n188), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n188), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n402), .B1(new_n425), .B2(new_n428), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n405), .B(KEYINPUT79), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n406), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(G469), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n320), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g264(.A(G113), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n453), .B2(new_n198), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n450), .A2(new_n454), .B1(new_n318), .B2(new_n319), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n383), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT85), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n449), .A2(KEYINPUT85), .A3(new_n456), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT6), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n449), .A2(new_n456), .A3(new_n458), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n449), .A2(KEYINPUT86), .A3(new_n456), .A4(new_n458), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n460), .A2(new_n457), .A3(new_n458), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n277), .A2(new_n215), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n215), .B1(new_n296), .B2(new_n303), .ZN(new_n473));
  OAI211_X1 g287(.A(G224), .B(new_n190), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n190), .A2(G224), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n471), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n477), .A2(KEYINPUT7), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n383), .B(new_n455), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n458), .B(KEYINPUT8), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n466), .A2(new_n467), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n491), .A3(new_n489), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n448), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT9), .B(G234), .ZN(new_n496));
  OAI21_X1  g310(.A(G221), .B1(new_n496), .B2(G902), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT78), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n446), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n452), .A2(G122), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n452), .A2(G122), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n370), .ZN(new_n504));
  XNOR2_X1  g318(.A(G128), .B(G143), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT13), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n270), .A2(G128), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(G134), .C1(KEYINPUT13), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n279), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT89), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n502), .B1(new_n501), .B2(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n370), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n505), .B(new_n279), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n503), .A2(new_n370), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n510), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n496), .A2(new_n187), .A3(G953), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n519), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n188), .ZN(new_n524));
  INV_X1    g338(.A(G478), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(KEYINPUT90), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(KEYINPUT90), .B2(new_n526), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n524), .B(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT17), .A3(G131), .ZN(new_n534));
  INV_X1    g348(.A(new_n532), .ZN(new_n535));
  OAI21_X1  g349(.A(G131), .B1(new_n535), .B2(new_n530), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n286), .A3(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n243), .A2(new_n238), .A3(new_n534), .A4(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n372), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT18), .A2(G131), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n531), .A2(new_n532), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n533), .A2(KEYINPUT18), .A3(G131), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n216), .A2(new_n218), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n223), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n544), .B(new_n545), .C1(new_n547), .C2(new_n234), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n540), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n542), .B1(new_n540), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n188), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G475), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n536), .A2(new_n537), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n233), .A2(KEYINPUT19), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n546), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n238), .B(new_n554), .C1(new_n557), .C2(G146), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n542), .B1(new_n558), .B2(new_n548), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n553), .B1(new_n549), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n548), .ZN(new_n561));
  INV_X1    g375(.A(new_n542), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n540), .A2(new_n542), .A3(new_n548), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT87), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G475), .A2(G902), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT20), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT88), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n529), .A2(new_n552), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G952), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G953), .ZN(new_n580));
  INV_X1    g394(.A(G234), .ZN(new_n581));
  INV_X1    g395(.A(G237), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT21), .B(G898), .Z(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT92), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n188), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n369), .A2(new_n500), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND3_X1  g406(.A1(new_n493), .A2(KEYINPUT93), .A3(new_n494), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n479), .A2(new_n489), .A3(new_n594), .A4(new_n491), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(new_n447), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n577), .A2(new_n552), .ZN(new_n598));
  AOI21_X1  g412(.A(G478), .B1(new_n522), .B2(new_n188), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT94), .B1(new_n519), .B2(new_n521), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(new_n522), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n525), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR4_X1   g419(.A1(new_n597), .A2(new_n589), .A3(new_n598), .A4(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n346), .B2(new_n188), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n335), .A2(new_n337), .ZN(new_n610));
  INV_X1    g424(.A(new_n345), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n342), .A2(KEYINPUT70), .A3(new_n343), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n348), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n262), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n499), .A3(new_n446), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n607), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n528), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n524), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n567), .B(KEYINPUT20), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n589), .B(KEYINPUT95), .Z(new_n624));
  AND4_X1   g438(.A1(new_n622), .A2(new_n623), .A3(new_n552), .A4(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n593), .A2(new_n625), .A3(new_n596), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n593), .A2(new_n625), .A3(new_n596), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT96), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n617), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(new_n193), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT36), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n245), .B(new_n634), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n260), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n255), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n500), .A2(new_n590), .A3(new_n615), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND2_X1  g454(.A1(new_n346), .A2(new_n349), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT32), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n346), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n368), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n425), .A2(new_n428), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n405), .B1(new_n646), .B2(new_n430), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n647), .B2(new_n429), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n439), .B1(new_n648), .B2(new_n437), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n498), .B1(new_n649), .B2(new_n445), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n584), .B1(new_n588), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n622), .A2(new_n623), .A3(new_n552), .A4(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n593), .A2(new_n654), .A3(new_n596), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n645), .A2(new_n650), .A3(new_n655), .A4(new_n637), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  INV_X1    g471(.A(new_n494), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n491), .B1(new_n479), .B2(new_n489), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n251), .A2(new_n189), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n248), .A2(new_n250), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT77), .A3(new_n253), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n663), .A2(new_n665), .B1(new_n260), .B2(new_n635), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n354), .A2(new_n343), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n362), .A2(new_n332), .A3(new_n343), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n188), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n643), .A2(new_n644), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n598), .A2(new_n448), .A3(new_n529), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n662), .A2(new_n666), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n652), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n650), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n650), .A2(KEYINPUT40), .A3(new_n674), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n270), .ZN(G45));
  NOR2_X1   g494(.A1(new_n598), .A2(new_n605), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n681), .A2(new_n593), .A3(new_n596), .A4(new_n653), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(new_n645), .A3(new_n650), .A4(new_n637), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  NAND2_X1  g498(.A1(new_n436), .A2(new_n188), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n497), .A3(new_n438), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n606), .A2(new_n369), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n629), .A2(new_n627), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n369), .A3(new_n688), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NOR2_X1   g508(.A1(new_n687), .A2(new_n597), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(new_n590), .A3(new_n645), .A4(new_n637), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n497), .A3(new_n438), .A4(new_n624), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n529), .B1(new_n552), .B2(new_n577), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n593), .A2(new_n596), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n363), .A2(new_n343), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n348), .B1(new_n610), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n609), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT97), .B1(new_n704), .B2(new_n616), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT97), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n609), .A2(new_n703), .A3(new_n262), .A4(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n701), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NOR3_X1   g523(.A1(new_n609), .A2(new_n666), .A3(new_n703), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n682), .A2(new_n710), .A3(new_n688), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(KEYINPUT98), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n384), .B1(new_n420), .B2(new_n421), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT12), .B1(new_n714), .B2(new_n397), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n401), .A2(new_n396), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n433), .B2(new_n434), .ZN(new_n718));
  INV_X1    g532(.A(new_n442), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n441), .A2(KEYINPUT98), .A3(new_n442), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(G469), .A3(new_n444), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n438), .A3(new_n440), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n658), .A2(new_n659), .A3(new_n448), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(new_n497), .A3(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n598), .A2(new_n605), .A3(new_n652), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR3_X1    g541(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT100), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT100), .B1(new_n350), .B2(new_n351), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n368), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n730), .A3(KEYINPUT42), .A4(new_n616), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n725), .A2(new_n645), .A3(new_n616), .A4(new_n726), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(KEYINPUT99), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT99), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  NAND3_X1  g551(.A1(new_n369), .A2(new_n654), .A3(new_n725), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G134), .ZN(G36));
  NAND2_X1  g553(.A1(new_n577), .A2(new_n552), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n605), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT43), .B1(new_n740), .B2(new_n605), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n637), .B1(new_n609), .B2(new_n614), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT102), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT102), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n637), .C1(new_n609), .C2(new_n614), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n724), .B1(new_n750), .B2(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n749), .ZN(new_n752));
  INV_X1    g566(.A(new_n745), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT44), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT103), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n750), .A2(new_n756), .A3(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n751), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n443), .A2(new_n444), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n437), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n444), .A4(new_n721), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n439), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n438), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n497), .B(new_n674), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND3_X1  g583(.A1(new_n726), .A2(new_n724), .A3(new_n262), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n645), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n497), .B(new_n774), .C1(new_n764), .C2(new_n765), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n497), .B1(new_n764), .B2(new_n765), .ZN(new_n776));
  INV_X1    g590(.A(new_n774), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n773), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n775), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n686), .A2(new_n438), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT107), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n498), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n584), .B(new_n753), .C1(new_n705), .C2(new_n707), .ZN(new_n786));
  INV_X1    g600(.A(new_n724), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(KEYINPUT112), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n778), .A2(new_n775), .B1(new_n498), .B2(new_n783), .ZN(new_n791));
  INV_X1    g605(.A(new_n788), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n743), .A2(new_n584), .A3(new_n744), .ZN(new_n794));
  INV_X1    g608(.A(new_n705), .ZN(new_n795));
  INV_X1    g609(.A(new_n707), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n660), .B(KEYINPUT38), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n448), .A3(new_n688), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT50), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n786), .B2(new_n799), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n688), .A2(new_n724), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n805), .A2(new_n583), .A3(new_n671), .A4(new_n262), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n598), .A2(new_n605), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n794), .A2(new_n687), .A3(new_n787), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n806), .A2(new_n808), .B1(new_n710), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n789), .A2(new_n793), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n812));
  AND2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n797), .B2(new_n800), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n786), .A2(new_n802), .A3(new_n799), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n785), .A2(new_n788), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n804), .A2(KEYINPUT113), .A3(new_n810), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(KEYINPUT51), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(new_n695), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n806), .A2(new_n681), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n580), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n730), .A2(new_n809), .A3(new_n616), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT48), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT48), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT114), .B1(new_n813), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n811), .A2(new_n812), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n821), .A4(new_n828), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n740), .A2(new_n605), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(new_n578), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n495), .A3(new_n624), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n615), .A2(new_n590), .A3(new_n637), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n446), .A2(new_n495), .A3(new_n499), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n617), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n500), .A2(new_n645), .A3(new_n590), .A4(new_n616), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT108), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n835), .A2(new_n495), .A3(new_n624), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n650), .A3(new_n616), .A4(new_n615), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT108), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n591), .A2(new_n843), .A3(new_n844), .A4(new_n638), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n689), .A2(new_n693), .A3(new_n708), .A4(new_n696), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n623), .A2(new_n529), .A3(new_n552), .A4(new_n653), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n787), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n650), .A3(new_n645), .A4(new_n637), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n725), .A2(new_n710), .A3(new_n726), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n738), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n736), .A2(new_n846), .A3(new_n847), .A4(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n593), .A2(new_n596), .A3(new_n699), .A4(new_n653), .ZN(new_n855));
  INV_X1    g669(.A(new_n497), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n649), .B2(new_n722), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n857), .A3(new_n671), .A4(new_n666), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n683), .A2(new_n656), .A3(new_n858), .A4(new_n711), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT52), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n732), .A2(new_n733), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n732), .A2(KEYINPUT99), .A3(new_n733), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n852), .B1(new_n869), .B2(new_n731), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n859), .A2(KEYINPUT109), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n859), .A2(KEYINPUT109), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n693), .A2(new_n708), .A3(new_n689), .A4(new_n696), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n845), .B2(new_n841), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n864), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n862), .B1(new_n854), .B2(new_n860), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n870), .A2(new_n875), .A3(KEYINPUT53), .A4(new_n877), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n830), .A2(new_n833), .A3(new_n882), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n579), .A2(new_n190), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT115), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n783), .B(KEYINPUT49), .Z(new_n891));
  NAND4_X1  g705(.A1(new_n616), .A2(new_n447), .A3(new_n499), .A4(new_n741), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT106), .Z(new_n893));
  OR4_X1    g707(.A1(new_n671), .A2(new_n891), .A3(new_n662), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n894), .ZN(G75));
  AOI21_X1  g709(.A(new_n188), .B1(new_n883), .B2(new_n885), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n470), .B(KEYINPUT116), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n478), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n897), .A2(new_n900), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n190), .A2(G952), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  NAND2_X1  g718(.A1(new_n883), .A2(new_n885), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n884), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n439), .B(KEYINPUT57), .Z(new_n907));
  OAI21_X1  g721(.A(new_n436), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n896), .A2(new_n762), .A3(new_n761), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND2_X1   g724(.A1(new_n560), .A2(new_n565), .ZN(new_n911));
  AND2_X1   g725(.A1(KEYINPUT58), .A2(G475), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n896), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n896), .B2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n903), .ZN(G60));
  NAND2_X1  g729(.A1(new_n882), .A2(new_n886), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n603), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n903), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n603), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n906), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT117), .Z(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n883), .B2(new_n885), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n259), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT119), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n928), .A2(new_n932), .A3(new_n259), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n920), .A2(KEYINPUT61), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n928), .A2(new_n936), .A3(new_n635), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n928), .B2(new_n635), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n920), .B1(new_n928), .B2(new_n259), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n905), .A2(new_n635), .A3(new_n926), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n928), .A2(new_n936), .A3(new_n635), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n934), .A2(new_n939), .B1(new_n944), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g759(.A(G224), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n587), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n877), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n898), .B1(G898), .B2(new_n190), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT120), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NAND2_X1  g765(.A1(new_n730), .A2(new_n616), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n700), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n767), .B1(new_n758), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n656), .A2(new_n711), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n683), .A3(new_n738), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n869), .B2(new_n731), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n954), .A2(new_n190), .A3(new_n779), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n313), .A2(new_n317), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT121), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n557), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n835), .B(KEYINPUT122), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n787), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n650), .A3(new_n369), .A4(new_n674), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n779), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n955), .A2(new_n683), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(new_n679), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n970), .A2(new_n679), .A3(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n969), .B(new_n768), .C1(new_n972), .C2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n190), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n964), .B(new_n965), .C1(new_n976), .C2(new_n961), .ZN(new_n977));
  INV_X1    g791(.A(new_n964), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n961), .B1(new_n975), .B2(new_n190), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT123), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n977), .B2(new_n981), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  INV_X1    g800(.A(new_n877), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n975), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n667), .ZN(new_n989));
  INV_X1    g803(.A(new_n881), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n355), .A2(new_n357), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n991), .A2(new_n992), .B1(new_n323), .B2(new_n334), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n986), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n989), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n954), .A2(new_n779), .A3(new_n877), .A4(new_n957), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n998), .A2(KEYINPUT124), .A3(new_n986), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT124), .B1(new_n998), .B2(new_n986), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n354), .A2(new_n343), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT125), .B1(new_n1002), .B2(new_n903), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1001), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n998), .A2(new_n986), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(KEYINPUT124), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1004), .B(new_n920), .C1(new_n1007), .C2(new_n999), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n997), .B1(new_n1003), .B2(new_n1008), .ZN(G57));
endmodule


