//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n463), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n475), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT68), .Z(G162));
  NAND2_X1  g063(.A1(new_n475), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n474), .A2(new_n463), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n463), .A2(new_n465), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n474), .A2(new_n463), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT69), .B(G51), .Z(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n510), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n511), .A2(new_n530), .B1(new_n513), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n511), .A2(new_n537), .B1(new_n513), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  AND2_X1   g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  NOR2_X1   g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n511), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT70), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT71), .B(G65), .Z(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n523), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n552), .A2(new_n557), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND3_X1  g139(.A1(new_n554), .A2(G87), .A3(new_n555), .ZN(new_n565));
  INV_X1    g140(.A(G74), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n508), .B1(new_n523), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(G49), .B2(new_n550), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G288));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  INV_X1    g145(.A(G73), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n549), .ZN(new_n572));
  NAND3_X1  g147(.A1(KEYINPUT72), .A2(G73), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n523), .C2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n550), .B2(G48), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n554), .A2(G86), .A3(new_n555), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT73), .Z(G305));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n523), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n508), .B1(new_n582), .B2(KEYINPUT74), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(KEYINPUT74), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n523), .A2(new_n548), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT75), .B(G85), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(new_n586), .B1(new_n550), .B2(G47), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G54), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n508), .B1(new_n591), .B2(new_n513), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n556), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(new_n540), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n597), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g187(.A1(new_n472), .A2(new_n463), .A3(new_n465), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n483), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n480), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n475), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT76), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT77), .Z(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT78), .Z(new_n643));
  NOR2_X1   g218(.A1(G2072), .A2(G2078), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n442), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(KEYINPUT17), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n641), .B(new_n642), .C1(new_n442), .C2(new_n644), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n647), .A3(new_n641), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT79), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n658), .A2(new_n663), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n659), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G25), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n483), .A2(G131), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n480), .A2(G119), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT81), .B1(G95), .B2(G2105), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g257(.A1(KEYINPUT81), .A2(G95), .A3(G2105), .ZN(new_n683));
  OAI221_X1 g258(.A(G2104), .B1(G107), .B2(new_n475), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n678), .B1(new_n686), .B2(new_n677), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  MUX2_X1   g264(.A(G24), .B(G290), .S(G16), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1986), .ZN(new_n691));
  AND2_X1   g266(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT82), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1971), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G23), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT84), .Z(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G288), .B2(new_n701), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n704), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n698), .B2(new_n699), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(KEYINPUT85), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n700), .A2(new_n716), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n694), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n715), .A2(KEYINPUT34), .A3(new_n717), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n701), .A2(G4), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n597), .B2(new_n701), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n483), .A2(G140), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n480), .A2(G128), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n475), .A2(G116), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n677), .A2(G26), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT87), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2067), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n701), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n540), .B2(new_n701), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(G1341), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n732), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  INV_X1    g326(.A(G127), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n493), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT89), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n483), .A2(G139), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G33), .B(new_n759), .S(G29), .Z(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2072), .Z(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n477), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2084), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  NOR2_X1   g343(.A1(new_n621), .A2(new_n677), .ZN(new_n769));
  INV_X1    g344(.A(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(KEYINPUT30), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n768), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n701), .A2(G21), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G168), .B2(new_n701), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n761), .A2(new_n767), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n701), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n701), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT91), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n677), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n677), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n781), .A2(new_n782), .B1(G2078), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT92), .B(G1956), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n701), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n601), .B2(new_n701), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n786), .B1(new_n782), .B2(new_n781), .C1(new_n787), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n677), .A2(G32), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G141), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n480), .A2(G129), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT26), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI22_X1  g374(.A1(G105), .A2(new_n472), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n794), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n793), .B1(new_n802), .B2(new_n677), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT27), .B(G1996), .Z(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT90), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n790), .A2(new_n787), .ZN(new_n807));
  INV_X1    g382(.A(G2078), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n784), .A2(new_n808), .B1(new_n803), .B2(new_n804), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n792), .A2(new_n806), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n748), .A2(new_n749), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n728), .A2(new_n750), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n724), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(G311));
  INV_X1    g390(.A(new_n814), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n816), .A2(new_n724), .A3(new_n812), .ZN(G150));
  NAND2_X1  g392(.A1(new_n597), .A2(G559), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT38), .Z(new_n819));
  AOI22_X1  g394(.A1(G93), .A2(new_n585), .B1(new_n550), .B2(G55), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT93), .B1(new_n821), .B2(new_n508), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n821), .A2(KEYINPUT93), .A3(new_n508), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(new_n606), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n540), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n819), .B(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n825), .A2(new_n832), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n621), .B(new_n477), .ZN(new_n838));
  XOR2_X1   g413(.A(G162), .B(new_n838), .Z(new_n839));
  AND3_X1   g414(.A1(new_n497), .A2(KEYINPUT94), .A3(new_n499), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT94), .B1(new_n497), .B2(new_n499), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n495), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n802), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n737), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n737), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(KEYINPUT4), .B2(new_n491), .ZN(new_n851));
  INV_X1    g426(.A(new_n841), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n497), .A2(KEYINPUT94), .A3(new_n499), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n849), .A2(new_n854), .A3(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n480), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n475), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G142), .B2(new_n483), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n614), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n685), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n848), .A2(new_n855), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n848), .B2(new_n855), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n839), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  INV_X1    g443(.A(new_n839), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n864), .B(new_n869), .C1(new_n866), .C2(KEYINPUT96), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n866), .A2(KEYINPUT96), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n867), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n829), .B(KEYINPUT97), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n610), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n609), .A2(new_n876), .A3(G299), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n878));
  NAND2_X1  g453(.A1(G299), .A2(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n597), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n877), .A2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n875), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(G305), .B(G166), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n893));
  XNOR2_X1  g468(.A(G290), .B(G288), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(KEYINPUT101), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n890), .A2(KEYINPUT42), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n891), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n891), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(G868), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n825), .ZN(G331));
  AND3_X1   g481(.A1(new_n827), .A2(G301), .A3(new_n828), .ZN(new_n907));
  AOI21_X1  g482(.A(G301), .B1(new_n827), .B2(new_n828), .ZN(new_n908));
  OAI21_X1  g483(.A(G286), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n829), .A2(G171), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n827), .A2(G301), .A3(new_n828), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(G168), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n888), .B2(new_n885), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n881), .B1(new_n909), .B2(new_n912), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n898), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n868), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n909), .A2(new_n912), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n889), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n899), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n916), .B2(new_n868), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n881), .A2(new_n884), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n883), .A2(new_n887), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n915), .B1(new_n928), .B2(KEYINPUT103), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n919), .A2(new_n930), .A3(new_n927), .A4(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n898), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n868), .A4(new_n921), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n925), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n899), .B1(new_n929), .B2(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n921), .A2(new_n868), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n937), .C2(new_n938), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n922), .A2(new_n923), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(KEYINPUT43), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n936), .B1(new_n944), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n842), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n468), .A2(G2105), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n472), .A2(G101), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(G40), .A3(new_n476), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n473), .A2(new_n954), .A3(G40), .A4(new_n476), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n737), .B(new_n743), .ZN(new_n958));
  INV_X1    g533(.A(G1996), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n801), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n686), .A2(new_n688), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n686), .A2(new_n688), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(G290), .B(G1986), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT123), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT109), .B(G8), .Z(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(G286), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n953), .A2(new_n955), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n842), .A2(new_n973), .A3(new_n946), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n946), .B1(new_n851), .B2(new_n500), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G2084), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n949), .A2(KEYINPUT111), .A3(new_n972), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n842), .B2(new_n946), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(new_n956), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n495), .B2(new_n501), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT45), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n985), .B2(new_n776), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n971), .B1(new_n987), .B2(new_n968), .ZN(new_n988));
  INV_X1    g563(.A(new_n984), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n956), .B1(new_n947), .B2(new_n948), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(KEYINPUT111), .ZN(new_n991));
  AOI21_X1  g566(.A(G1966), .B1(new_n991), .B2(new_n982), .ZN(new_n992));
  OAI21_X1  g567(.A(G8), .B1(new_n992), .B2(new_n978), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n970), .B1(new_n993), .B2(new_n969), .ZN(new_n994));
  OAI211_X1 g569(.A(G286), .B(new_n968), .C1(new_n992), .C2(new_n978), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n988), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n998));
  INV_X1    g573(.A(G1971), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n953), .B(new_n955), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT106), .B(G2090), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n972), .A2(new_n974), .A3(new_n976), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  NAND4_X1  g585(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AND4_X1   g587(.A1(new_n998), .A2(new_n1005), .A3(G8), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n998), .B1(new_n1015), .B2(new_n1012), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n842), .A2(new_n953), .A3(new_n946), .A4(new_n955), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n565), .A2(new_n568), .A3(G1976), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n968), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(KEYINPUT110), .A3(new_n968), .A4(new_n1019), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(KEYINPUT52), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n576), .A2(new_n577), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n572), .A2(new_n573), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n574), .B1(new_n504), .B2(new_n505), .ZN(new_n1028));
  OAI21_X1  g603(.A(G651), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n550), .A2(G48), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n506), .A2(new_n510), .A3(G86), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G1981), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1026), .A2(new_n1033), .A3(KEYINPUT49), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n968), .A3(new_n1018), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1018), .A2(new_n968), .A3(new_n1019), .A4(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n973), .B(new_n946), .C1(new_n851), .C2(new_n500), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1043), .A2(new_n953), .A3(new_n955), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1003), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n967), .B1(new_n1002), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1024), .B(new_n1042), .C1(new_n1047), .C2(new_n1012), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n997), .B1(new_n1017), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT45), .B1(new_n502), .B2(new_n946), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n956), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AND4_X1   g628(.A1(new_n974), .A2(new_n972), .A3(new_n976), .A4(new_n1003), .ZN(new_n1054));
  OAI211_X1 g629(.A(G8), .B(new_n1012), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT108), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1015), .A2(new_n998), .A3(new_n1012), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1024), .A2(new_n1042), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1002), .A2(new_n1046), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1012), .B1(new_n1060), .B2(new_n968), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1062), .A3(KEYINPUT120), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n975), .A2(new_n948), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n972), .A2(new_n1052), .A3(new_n808), .A4(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT117), .B(G1961), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1066), .A2(new_n1067), .B1(new_n977), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT119), .B(G2078), .Z(new_n1071));
  NOR3_X1   g646(.A1(new_n952), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n949), .A2(new_n1052), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1070), .A2(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n979), .A2(new_n982), .A3(new_n984), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1064), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n996), .A2(new_n1049), .A3(new_n1063), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1064), .B1(new_n1074), .B2(G171), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1069), .A2(new_n1077), .A3(G301), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT121), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1069), .A2(new_n1077), .A3(new_n1084), .A4(G301), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT122), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n966), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1049), .A2(new_n1063), .A3(new_n1079), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1086), .B(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1089), .A2(new_n1091), .A3(KEYINPUT123), .A4(new_n996), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT112), .B(G1956), .Z(new_n1096));
  AOI22_X1  g671(.A1(new_n1093), .A2(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n552), .B2(KEYINPUT113), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(G299), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1018), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n977), .A2(new_n731), .B1(new_n1102), .B2(new_n743), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n609), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT114), .Z(new_n1106));
  INV_X1    g681(.A(new_n1100), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1107), .A2(new_n1101), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1107), .B2(new_n1101), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n597), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1109), .B(new_n1110), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT115), .B(G1996), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT58), .B(G1341), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1102), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(KEYINPUT116), .A3(new_n540), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT59), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n597), .B2(new_n1112), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1106), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1088), .A2(new_n1092), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n969), .B1(new_n986), .B2(new_n1014), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n995), .A3(KEYINPUT51), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n970), .B(new_n969), .C1(new_n986), .C2(new_n967), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1058), .A2(KEYINPUT120), .A3(new_n1062), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(new_n1132), .A3(KEYINPUT124), .A4(new_n1078), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1049), .A2(new_n1063), .A3(new_n1078), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT62), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1038), .A2(new_n1039), .A3(new_n565), .A4(new_n568), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n967), .B(new_n1102), .C1(new_n1140), .C2(new_n1026), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1061), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n986), .A2(new_n967), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1059), .B1(new_n1144), .B2(new_n1058), .ZN(new_n1145));
  OAI21_X1  g720(.A(G168), .B1(new_n1015), .B2(new_n1012), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1059), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1143), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1141), .B(new_n1145), .C1(KEYINPUT63), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n965), .B1(new_n1123), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n963), .A2(new_n957), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT126), .Z(new_n1153));
  NOR4_X1   g728(.A1(new_n949), .A2(G1986), .A3(new_n956), .A4(G290), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n958), .A2(new_n802), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n957), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT125), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n957), .A2(new_n959), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT46), .Z(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n958), .A2(new_n960), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1164), .A2(new_n961), .B1(G2067), .B2(new_n737), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1156), .B(new_n1163), .C1(new_n957), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1151), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g742(.A1(G227), .A2(new_n460), .ZN(new_n1169));
  AND2_X1   g743(.A1(new_n639), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g744(.A1(new_n1170), .A2(KEYINPUT127), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT127), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n675), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n924), .A2(new_n935), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n1173), .A2(new_n872), .A3(new_n1174), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


