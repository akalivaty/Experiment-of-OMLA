

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(n390), .B(n389), .ZN(n392) );
  XNOR2_X1 U324 ( .A(KEYINPUT119), .B(n449), .ZN(n556) );
  XOR2_X1 U325 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n291) );
  XNOR2_X1 U326 ( .A(n388), .B(KEYINPUT73), .ZN(n389) );
  NOR2_X1 U327 ( .A1(n464), .A2(n561), .ZN(n447) );
  XNOR2_X1 U328 ( .A(n424), .B(n423), .ZN(n446) );
  XNOR2_X1 U329 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U330 ( .A(n399), .B(n398), .ZN(n569) );
  INV_X1 U331 ( .A(G183GAT), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n450), .B(KEYINPUT120), .ZN(n451) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT81), .B(G64GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G211GAT), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U337 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT80), .B(KEYINPUT12), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U341 ( .A(G22GAT), .B(G155GAT), .Z(n335) );
  XOR2_X1 U342 ( .A(n335), .B(G71GAT), .Z(n299) );
  XOR2_X1 U343 ( .A(G1GAT), .B(G8GAT), .Z(n367) );
  XNOR2_X1 U344 ( .A(n367), .B(G183GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n304) );
  XNOR2_X1 U346 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n300), .B(KEYINPUT72), .ZN(n391) );
  XOR2_X1 U348 ( .A(n391), .B(KEYINPUT15), .Z(n302) );
  NAND2_X1 U349 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n306) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n575) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n310) );
  XNOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U358 ( .A(n311), .B(G183GAT), .Z(n313) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(G176GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n413) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G71GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n314), .B(G120GAT), .ZN(n385) );
  XOR2_X1 U363 ( .A(KEYINPUT20), .B(n385), .Z(n316) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n319) );
  XNOR2_X1 U366 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n317) );
  XOR2_X1 U367 ( .A(KEYINPUT0), .B(G127GAT), .Z(n439) );
  XNOR2_X1 U368 ( .A(n317), .B(n439), .ZN(n318) );
  XOR2_X1 U369 ( .A(n319), .B(n318), .Z(n321) );
  XOR2_X1 U370 ( .A(G113GAT), .B(G15GAT), .Z(n370) );
  XOR2_X1 U371 ( .A(G43GAT), .B(G134GAT), .Z(n350) );
  XNOR2_X1 U372 ( .A(n370), .B(n350), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X2 U374 ( .A(n413), .B(n322), .ZN(n525) );
  XNOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n323), .B(KEYINPUT21), .ZN(n324) );
  XOR2_X1 U377 ( .A(n324), .B(KEYINPUT89), .Z(n326) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n412) );
  XOR2_X1 U380 ( .A(G50GAT), .B(G162GAT), .Z(n356) );
  XOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT91), .Z(n328) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n438) );
  XOR2_X1 U384 ( .A(n356), .B(n438), .Z(n330) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n412), .B(n331), .ZN(n343) );
  XOR2_X1 U388 ( .A(KEYINPUT93), .B(KEYINPUT87), .Z(n333) );
  XNOR2_X1 U389 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U391 ( .A(n334), .B(KEYINPUT92), .Z(n337) );
  XNOR2_X1 U392 ( .A(n335), .B(KEYINPUT24), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U394 ( .A(n338), .B(G204GAT), .Z(n341) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(G78GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n339), .B(G148GAT), .ZN(n384) );
  XNOR2_X1 U397 ( .A(n384), .B(KEYINPUT22), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n464) );
  XNOR2_X1 U400 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n411) );
  XOR2_X1 U401 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n345) );
  XNOR2_X1 U402 ( .A(G218GAT), .B(KEYINPUT76), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U404 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U407 ( .A(n349), .B(n348), .Z(n352) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G92GAT), .Z(n393) );
  XNOR2_X1 U409 ( .A(n350), .B(n393), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U411 ( .A(G36GAT), .B(KEYINPUT79), .Z(n416) );
  XOR2_X1 U412 ( .A(n353), .B(n416), .Z(n358) );
  XOR2_X1 U413 ( .A(G29GAT), .B(KEYINPUT8), .Z(n355) );
  XNOR2_X1 U414 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n371) );
  XNOR2_X1 U416 ( .A(n371), .B(n356), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U418 ( .A(G106GAT), .B(G99GAT), .Z(n360) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(G190GAT), .B(n361), .Z(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n534) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G141GAT), .Z(n365) );
  XNOR2_X1 U424 ( .A(G50GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U426 ( .A(n366), .B(G43GAT), .Z(n369) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(n367), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U429 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U433 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n377) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U436 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n379) );
  XNOR2_X1 U437 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n563) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n390) );
  XNOR2_X1 U442 ( .A(KEYINPUT33), .B(KEYINPUT75), .ZN(n387) );
  AND2_X1 U443 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n392), .B(n391), .ZN(n399) );
  XOR2_X1 U446 ( .A(G204GAT), .B(G64GAT), .Z(n418) );
  XNOR2_X1 U447 ( .A(n393), .B(n418), .ZN(n397) );
  XOR2_X1 U448 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n395) );
  XNOR2_X1 U449 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT41), .B(n569), .ZN(n552) );
  NOR2_X1 U452 ( .A1(n563), .A2(n552), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n400), .B(n291), .ZN(n401) );
  NAND2_X1 U454 ( .A1(n401), .A2(n575), .ZN(n402) );
  NOR2_X1 U455 ( .A1(n534), .A2(n402), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n403), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n404), .B(n534), .ZN(n580) );
  NOR2_X1 U459 ( .A1(n575), .A2(n580), .ZN(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT45), .B(n405), .Z(n406) );
  NOR2_X1 U461 ( .A1(n569), .A2(n406), .ZN(n407) );
  NAND2_X1 U462 ( .A1(n407), .A2(n563), .ZN(n408) );
  NAND2_X1 U463 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n521) );
  XNOR2_X1 U465 ( .A(n413), .B(n412), .ZN(n422) );
  XOR2_X1 U466 ( .A(G92GAT), .B(KEYINPUT97), .Z(n415) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U470 ( .A(G8GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U472 ( .A(n422), .B(n421), .ZN(n455) );
  NAND2_X1 U473 ( .A1(n521), .A2(n455), .ZN(n424) );
  XOR2_X1 U474 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n423) );
  XOR2_X1 U475 ( .A(G85GAT), .B(G120GAT), .Z(n426) );
  XNOR2_X1 U476 ( .A(G113GAT), .B(G134GAT), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(G155GAT), .Z(n428) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U481 ( .A(n430), .B(n429), .Z(n435) );
  XOR2_X1 U482 ( .A(KEYINPUT6), .B(G57GAT), .Z(n432) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(KEYINPUT1), .B(n433), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n445) );
  XOR2_X1 U487 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n437) );
  XNOR2_X1 U488 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U490 ( .A(n438), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U491 ( .A(G29GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U493 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X1 U494 ( .A(n445), .B(n444), .ZN(n510) );
  NAND2_X1 U495 ( .A1(n446), .A2(n510), .ZN(n561) );
  XNOR2_X1 U496 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NOR2_X1 U497 ( .A1(n525), .A2(n448), .ZN(n449) );
  NOR2_X1 U498 ( .A1(n575), .A2(n556), .ZN(n452) );
  NOR2_X1 U499 ( .A1(n563), .A2(n569), .ZN(n485) );
  XOR2_X1 U500 ( .A(n455), .B(KEYINPUT27), .Z(n465) );
  XOR2_X1 U501 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n454) );
  NAND2_X1 U502 ( .A1(n464), .A2(n525), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(n562) );
  NOR2_X1 U504 ( .A1(n465), .A2(n562), .ZN(n460) );
  INV_X1 U505 ( .A(n455), .ZN(n513) );
  NOR2_X1 U506 ( .A1(n525), .A2(n513), .ZN(n456) );
  NOR2_X1 U507 ( .A1(n464), .A2(n456), .ZN(n457) );
  XOR2_X1 U508 ( .A(n457), .B(KEYINPUT100), .Z(n458) );
  XNOR2_X1 U509 ( .A(KEYINPUT25), .B(n458), .ZN(n459) );
  NOR2_X1 U510 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n461), .B(KEYINPUT101), .ZN(n462) );
  NAND2_X1 U512 ( .A1(n462), .A2(n510), .ZN(n463) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(n463), .Z(n470) );
  XNOR2_X1 U514 ( .A(n464), .B(KEYINPUT28), .ZN(n479) );
  XNOR2_X1 U515 ( .A(KEYINPUT86), .B(n525), .ZN(n466) );
  NOR2_X1 U516 ( .A1(n465), .A2(n510), .ZN(n520) );
  NAND2_X1 U517 ( .A1(n466), .A2(n520), .ZN(n467) );
  NOR2_X1 U518 ( .A1(n479), .A2(n467), .ZN(n468) );
  XNOR2_X1 U519 ( .A(n468), .B(KEYINPUT98), .ZN(n469) );
  NOR2_X1 U520 ( .A1(n470), .A2(n469), .ZN(n482) );
  XOR2_X1 U521 ( .A(KEYINPUT83), .B(KEYINPUT16), .Z(n472) );
  INV_X1 U522 ( .A(n534), .ZN(n557) );
  INV_X1 U523 ( .A(n575), .ZN(n531) );
  NAND2_X1 U524 ( .A1(n557), .A2(n531), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U526 ( .A1(n482), .A2(n473), .ZN(n498) );
  NAND2_X1 U527 ( .A1(n485), .A2(n498), .ZN(n480) );
  NOR2_X1 U528 ( .A1(n510), .A2(n480), .ZN(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(n474), .Z(n475) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U531 ( .A1(n513), .A2(n480), .ZN(n476) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n525), .A2(n480), .ZN(n478) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  INV_X1 U536 ( .A(n479), .ZN(n523) );
  NOR2_X1 U537 ( .A1(n523), .A2(n480), .ZN(n481) );
  XOR2_X1 U538 ( .A(G22GAT), .B(n481), .Z(G1327GAT) );
  NOR2_X1 U539 ( .A1(n482), .A2(n580), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n575), .A2(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n484), .ZN(n509) );
  NAND2_X1 U542 ( .A1(n509), .A2(n485), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT38), .B(n486), .ZN(n494) );
  NOR2_X1 U544 ( .A1(n510), .A2(n494), .ZN(n490) );
  XOR2_X1 U545 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n488) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT104), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n494), .A2(n513), .ZN(n491) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n525), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(n492), .Z(n493) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n523), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  INV_X1 U558 ( .A(n563), .ZN(n526) );
  NOR2_X1 U559 ( .A1(n552), .A2(n526), .ZN(n508) );
  NAND2_X1 U560 ( .A1(n508), .A2(n498), .ZN(n505) );
  NOR2_X1 U561 ( .A1(n510), .A2(n505), .ZN(n499) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n513), .A2(n505), .ZN(n502) );
  XNOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U567 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  NOR2_X1 U568 ( .A1(n525), .A2(n505), .ZN(n504) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n523), .A2(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n510), .A2(n516), .ZN(n511) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT110), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n516), .ZN(n514) );
  XOR2_X1 U578 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U579 ( .A1(n525), .A2(n516), .ZN(n515) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U581 ( .A1(n523), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT113), .ZN(n540) );
  NAND2_X1 U587 ( .A1(n523), .A2(n540), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  INV_X1 U592 ( .A(n552), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n535), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n535), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n537) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  INV_X1 U602 ( .A(n562), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n563), .A2(n548), .ZN(n541) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  NOR2_X1 U606 ( .A1(n548), .A2(n552), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n575), .A2(n548), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(n546), .Z(n547) );
  XNOR2_X1 U613 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n557), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G162GAT), .B(KEYINPUT117), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n563), .A2(n556), .ZN(n551) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n551), .Z(G1348GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n556), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  OR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n579) );
  NOR2_X1 U628 ( .A1(n563), .A2(n579), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT59), .B(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  INV_X1 U634 ( .A(n569), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n579), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

