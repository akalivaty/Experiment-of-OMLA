//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n203), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(new_n203), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n209), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n211), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n233), .B(new_n236), .C1(new_n224), .C2(new_n225), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n227), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n202), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT67), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G97), .B(G107), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NAND3_X1  g0054(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n231), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n208), .A2(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G50), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n209), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n209), .A2(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(G20), .B2(new_n204), .ZN(new_n268));
  INV_X1    g0068(.A(new_n258), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n261), .B1(G50), .B2(new_n255), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT69), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(new_n276), .B2(new_n279), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT68), .B(G226), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(KEYINPUT70), .B(new_n277), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G222), .A2(G1698), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G223), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n294), .C1(G77), .C2(new_n289), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n287), .A2(new_n288), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n271), .B(new_n297), .C1(new_n298), .C2(new_n296), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n296), .A2(G179), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n270), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n259), .ZN(new_n307));
  INV_X1    g0107(.A(new_n262), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n260), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n307), .A2(new_n309), .B1(new_n255), .B2(new_n308), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT72), .A3(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT72), .B1(new_n312), .B2(G33), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n311), .B(new_n209), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G68), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n313), .A3(new_n314), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n321), .B2(new_n209), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT73), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n320), .A2(new_n313), .A3(new_n314), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT7), .B1(new_n324), .B2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(G68), .A4(new_n317), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G58), .A2(G68), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n209), .B1(new_n228), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G159), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n266), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n329), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n323), .A2(new_n327), .A3(KEYINPUT16), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n312), .A2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n314), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n339), .B2(new_n209), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n311), .B(G20), .C1(new_n338), .C2(new_n314), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n332), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n269), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n310), .B1(new_n337), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  OR2_X1    g0147(.A1(G223), .A2(G1698), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G226), .B2(new_n291), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n321), .A2(new_n349), .B1(new_n265), .B2(new_n214), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n294), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n276), .A2(new_n279), .ZN(new_n352));
  INV_X1    g0152(.A(G232), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G190), .B2(new_n357), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n346), .A2(new_n347), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n347), .B1(new_n346), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT17), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n337), .A2(new_n345), .ZN(new_n365));
  INV_X1    g0165(.A(new_n310), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n302), .B1(new_n351), .B2(new_n356), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n364), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n346), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT17), .B1(new_n346), .B2(new_n360), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n363), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n256), .A2(new_n203), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT12), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n203), .A2(G20), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n382), .B1(new_n263), .B2(new_n218), .C1(new_n201), .C2(new_n266), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n259), .A2(G68), .A3(new_n260), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT11), .B1(new_n383), .B2(new_n258), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT14), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G226), .A2(G1698), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n353), .B2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n392), .B1(new_n394), .B2(new_n289), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n277), .B1(new_n395), .B2(new_n276), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n352), .A2(KEYINPUT69), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n213), .B1(new_n397), .B2(new_n280), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n396), .A2(new_n398), .A3(KEYINPUT13), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n353), .A2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G226), .B2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n391), .B1(new_n402), .B2(new_n339), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n355), .B1(new_n403), .B2(new_n294), .ZN(new_n404));
  OAI21_X1  g0204(.A(G238), .B1(new_n281), .B2(new_n282), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n390), .B(G169), .C1(new_n399), .C2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT13), .B1(new_n396), .B2(new_n398), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(G179), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n409), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n390), .B1(new_n412), .B2(G169), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n389), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n289), .A2(G232), .A3(new_n291), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n220), .B2(new_n289), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n339), .A2(new_n213), .A3(new_n291), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n294), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n277), .C1(new_n219), .C2(new_n283), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n302), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT71), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n256), .A2(new_n218), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G20), .A2(G77), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n425), .B1(new_n262), .B2(new_n266), .C1(new_n263), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n258), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n419), .A2(G179), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n412), .A2(G200), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n388), .C1(new_n298), .C2(new_n412), .ZN(new_n434));
  INV_X1    g0234(.A(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n419), .A2(G200), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n436), .C1(new_n298), .C2(new_n419), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n414), .A2(new_n432), .A3(new_n434), .A4(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n306), .A2(new_n379), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n208), .A2(G45), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT5), .A2(G41), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n294), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n276), .A2(G274), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n445), .A2(G270), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n221), .A2(G1698), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G257), .B2(G1698), .ZN(new_n451));
  INV_X1    g0251(.A(G303), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n321), .A2(new_n451), .B1(new_n452), .B2(new_n289), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n294), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n256), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n208), .A2(G33), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n255), .A2(new_n458), .A3(new_n231), .A4(new_n257), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n456), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n257), .A2(new_n231), .B1(G20), .B2(new_n456), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n209), .C1(G33), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(KEYINPUT20), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n464), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n455), .A2(new_n470), .A3(KEYINPUT80), .A4(G179), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n449), .A2(new_n454), .A3(G179), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n469), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n449), .A2(new_n454), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(new_n469), .C1(new_n298), .C2(new_n476), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n470), .A2(new_n476), .A3(KEYINPUT21), .A4(G169), .ZN(new_n482));
  AND4_X1   g0282(.A1(new_n475), .A2(new_n478), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n445), .A2(G257), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n447), .A2(new_n448), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n219), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT4), .B1(new_n324), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n338), .A2(new_n314), .A3(G250), .A4(G1698), .ZN(new_n490));
  AND2_X1   g0290(.A1(KEYINPUT4), .A2(G244), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n338), .A2(new_n314), .A3(new_n491), .A4(new_n291), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n492), .A3(new_n462), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n294), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT77), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n490), .A2(new_n492), .A3(new_n462), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  INV_X1    g0298(.A(new_n488), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n321), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n276), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(KEYINPUT77), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n487), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n463), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n209), .B1(new_n218), .B2(new_n266), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n311), .B1(new_n289), .B2(G20), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n220), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n258), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n459), .A2(KEYINPUT76), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n459), .A2(KEYINPUT76), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(G97), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n256), .A2(new_n463), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n501), .A2(new_n486), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(G190), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n302), .B1(new_n501), .B2(new_n486), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n368), .B(new_n487), .C1(new_n496), .C2(new_n502), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n504), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n215), .A2(new_n291), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G257), .B2(new_n291), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n321), .A2(new_n526), .B1(new_n265), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n294), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n445), .A2(G264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n485), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n358), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n528), .A2(new_n294), .B1(new_n445), .B2(G264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n298), .A3(new_n485), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n514), .A2(G107), .A3(new_n515), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n255), .A2(G107), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT25), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n214), .A2(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n338), .A3(new_n314), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n209), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AND2_X1   g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(new_n209), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n320), .A2(new_n313), .A3(new_n209), .A4(new_n314), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n542), .A2(new_n214), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT24), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n313), .A2(new_n314), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(new_n209), .A3(new_n320), .A4(new_n551), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n543), .A4(new_n548), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n539), .B1(new_n559), .B2(new_n258), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n535), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n531), .A2(new_n302), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n533), .A2(new_n368), .A3(new_n485), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n269), .B1(new_n554), .B2(new_n558), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n539), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g0366(.A1(KEYINPUT78), .A2(G87), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT78), .A2(G87), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n391), .B2(new_n209), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n263), .B2(new_n463), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n203), .C2(new_n550), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n258), .B1(new_n256), .B2(new_n426), .ZN(new_n576));
  INV_X1    g0376(.A(new_n426), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n514), .A2(new_n577), .A3(new_n515), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n219), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G238), .B2(G1698), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n321), .A2(new_n581), .B1(new_n265), .B2(new_n456), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n294), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n276), .A2(G250), .A3(new_n440), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n446), .B2(new_n440), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n302), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n582), .B2(new_n294), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n368), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n579), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT79), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n589), .A2(new_n592), .A3(G190), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n589), .B2(G190), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n514), .A2(G87), .A3(new_n515), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n576), .B(new_n596), .C1(new_n358), .C2(new_n589), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n566), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n439), .A2(new_n483), .A3(new_n524), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT81), .ZN(G372));
  NOR2_X1   g0401(.A1(new_n589), .A2(new_n358), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n575), .A2(new_n258), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n426), .A2(new_n256), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n596), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n576), .A2(KEYINPUT82), .A3(new_n596), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT83), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n609), .A2(new_n610), .B1(new_n593), .B2(new_n594), .ZN(new_n611));
  AOI211_X1 g0411(.A(KEYINPUT83), .B(new_n602), .C1(new_n607), .C2(new_n608), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n475), .A2(new_n565), .A3(new_n481), .A4(new_n482), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n522), .A2(new_n523), .ZN(new_n615));
  INV_X1    g0415(.A(new_n518), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n519), .A2(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n494), .A2(new_n495), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n501), .A2(KEYINPUT77), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n486), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n616), .B(new_n617), .C1(new_n620), .C2(new_n358), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n614), .A2(new_n615), .A3(new_n621), .A4(new_n561), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n591), .B1(new_n613), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n615), .A2(new_n598), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n522), .A2(new_n523), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n626), .B(new_n591), .C1(new_n611), .C2(new_n612), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n627), .B2(new_n624), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n439), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g0429(.A(new_n629), .B(KEYINPUT84), .Z(new_n630));
  INV_X1    g0430(.A(new_n304), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n365), .A2(new_n360), .A3(new_n366), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT75), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n346), .A2(new_n347), .A3(new_n360), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n376), .B1(new_n635), .B2(KEYINPUT17), .ZN(new_n636));
  INV_X1    g0436(.A(new_n434), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n414), .B1(new_n432), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n373), .B2(new_n374), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n367), .A2(new_n364), .A3(new_n372), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT18), .B1(new_n346), .B2(new_n371), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(KEYINPUT85), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n631), .B1(new_n646), .B2(new_n300), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n630), .A2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n469), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n483), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n654), .B1(new_n564), .B2(new_n539), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n561), .A2(new_n565), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT87), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n561), .A2(new_n667), .A3(new_n565), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n565), .A2(new_n655), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n669), .A2(KEYINPUT88), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n663), .A2(G330), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n565), .A2(new_n654), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n659), .A2(new_n655), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n678), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n234), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n570), .A2(G116), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G1), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n229), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n655), .B1(new_n628), .B2(new_n623), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT90), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT90), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n693), .B(new_n655), .C1(new_n628), .C2(new_n623), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n615), .A2(new_n598), .A3(KEYINPUT26), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n697), .B(new_n591), .C1(new_n613), .C2(new_n622), .ZN(new_n698));
  OAI211_X1 g0498(.A(KEYINPUT29), .B(new_n655), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n599), .A2(new_n524), .A3(new_n483), .A4(new_n655), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n473), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n533), .A2(new_n589), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n449), .A2(new_n454), .A3(KEYINPUT89), .A4(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n704), .A3(new_n519), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n519), .A2(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n531), .A2(new_n476), .A3(new_n587), .A4(new_n368), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n709), .A2(new_n710), .B1(new_n620), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n654), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT31), .B(new_n654), .C1(new_n708), .C2(new_n712), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n701), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n700), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n689), .B1(new_n720), .B2(G1), .ZN(G364));
  INV_X1    g0521(.A(G13), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G45), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n684), .A2(new_n725), .A3(new_n208), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n265), .A3(KEYINPUT93), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT93), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G13), .B2(G33), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n231), .B1(G20), .B2(new_n302), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n250), .A2(G45), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT92), .Z(new_n736));
  NOR2_X1   g0536(.A1(new_n683), .A2(new_n324), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(G45), .C2(new_n229), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n683), .A2(new_n339), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n739), .A2(G355), .B1(new_n456), .B2(new_n683), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n733), .B(new_n734), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n209), .A2(G190), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT95), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(G159), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n749), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n747), .B2(new_n330), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(new_n368), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(G190), .A3(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n750), .B(new_n752), .C1(new_n201), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n368), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n742), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n760), .A2(G20), .A3(G190), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n289), .B1(new_n761), .B2(new_n218), .C1(new_n202), .C2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n753), .A2(new_n298), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n209), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n298), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n203), .B1(new_n766), .B2(new_n220), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n209), .B1(new_n743), .B2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n463), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n567), .B2(new_n569), .ZN(new_n771));
  OR4_X1    g0571(.A1(new_n763), .A2(new_n767), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n748), .A2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(new_n764), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT33), .B(G317), .ZN(new_n775));
  INV_X1    g0575(.A(new_n770), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(G303), .ZN(new_n777));
  INV_X1    g0577(.A(new_n766), .ZN(new_n778));
  INV_X1    g0578(.A(new_n768), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n778), .A2(G283), .B1(new_n779), .B2(G294), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n339), .B1(new_n762), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n761), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G311), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n773), .A2(new_n777), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n758), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n759), .A2(new_n772), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n727), .B(new_n741), .C1(new_n734), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n733), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n661), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n726), .B1(new_n663), .B2(G330), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G330), .B2(new_n663), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  AND4_X1   g0595(.A1(new_n429), .A2(new_n431), .A3(new_n420), .A4(new_n655), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n437), .B1(new_n435), .B2(new_n655), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(new_n797), .B2(new_n432), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n691), .A2(new_n694), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n655), .B(new_n798), .C1(new_n628), .C2(new_n623), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n726), .B1(new_n802), .B2(new_n718), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n718), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n731), .A2(new_n734), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n726), .B1(G77), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT97), .Z(new_n808));
  INV_X1    g0608(.A(new_n734), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n769), .B1(G283), .B2(new_n774), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n214), .B2(new_n766), .C1(new_n220), .C2(new_n770), .ZN(new_n811));
  INV_X1    g0611(.A(new_n762), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n289), .B1(new_n812), .B2(G294), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n456), .B2(new_n761), .C1(new_n747), .C2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n811), .B(new_n815), .C1(G303), .C2(new_n786), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n812), .A2(G143), .B1(new_n783), .B2(G159), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n264), .B2(new_n764), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G137), .B2(new_n786), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n321), .B1(new_n776), .B2(G50), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n766), .A2(new_n203), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G58), .B2(new_n779), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n821), .B(new_n823), .C1(new_n747), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n819), .B2(KEYINPUT34), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n816), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n808), .B1(new_n809), .B2(new_n827), .C1(new_n798), .C2(new_n732), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n804), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT98), .ZN(G384));
  INV_X1    g0630(.A(new_n508), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT35), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT35), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n832), .A2(G116), .A3(new_n232), .A4(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT36), .Z(new_n835));
  NAND3_X1  g0635(.A1(new_n230), .A2(G77), .A3(new_n328), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n201), .A2(G68), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n208), .B(G13), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT39), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n641), .A2(new_n363), .A3(new_n377), .A4(new_n644), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n346), .A2(new_n652), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n367), .A2(new_n372), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n632), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n845), .B2(new_n842), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT37), .B1(new_n367), .B2(new_n372), .ZN(new_n847));
  INV_X1    g0647(.A(new_n842), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(new_n633), .A3(new_n634), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT38), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n323), .A2(new_n327), .A3(new_n336), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(KEYINPUT100), .A3(new_n344), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n344), .A2(KEYINPUT100), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n323), .A2(new_n327), .A3(new_n336), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n853), .A2(new_n258), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n652), .B1(new_n856), .B2(new_n366), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n378), .A2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n856), .A2(new_n366), .B1(new_n371), .B2(new_n652), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n635), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n849), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n840), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n414), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n655), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n858), .A2(new_n861), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n863), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n652), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n645), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(new_n870), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n389), .A2(new_n654), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n414), .A2(KEYINPUT99), .A3(new_n434), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT99), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n414), .A2(new_n878), .A3(new_n434), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n411), .A2(new_n876), .A3(new_n413), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n876), .A2(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n796), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n801), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n874), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n872), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n695), .A2(new_n439), .A3(new_n699), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n647), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n886), .B(new_n888), .Z(new_n889));
  AND3_X1   g0689(.A1(new_n701), .A2(new_n715), .A3(new_n716), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n877), .A2(new_n876), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n879), .A2(new_n880), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n798), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n858), .B2(new_n861), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n862), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n841), .A2(new_n842), .B1(new_n849), .B2(new_n846), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n870), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n890), .B2(new_n893), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n717), .A2(new_n881), .A3(KEYINPUT101), .A4(new_n798), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n439), .A2(new_n717), .ZN(new_n906));
  OAI21_X1  g0706(.A(G330), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n889), .A2(new_n908), .B1(new_n208), .B2(new_n723), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n889), .A2(new_n908), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n839), .B1(new_n909), .B2(new_n910), .ZN(G367));
  NAND3_X1  g0711(.A1(new_n607), .A2(new_n608), .A3(new_n654), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n591), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT102), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n591), .B(new_n912), .C1(new_n611), .C2(new_n612), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n733), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n733), .A2(new_n734), .ZN(new_n919));
  INV_X1    g0719(.A(new_n737), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n919), .B1(new_n234), .B2(new_n426), .C1(new_n920), .C2(new_n245), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n726), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT107), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n774), .A2(G159), .B1(new_n783), .B2(G50), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n786), .A2(G143), .B1(KEYINPUT108), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n748), .A2(G137), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n289), .B1(new_n762), .B2(new_n264), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n202), .A2(new_n770), .B1(new_n766), .B2(new_n218), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(G68), .C2(new_n779), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n927), .A2(new_n928), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G283), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n321), .B1(new_n761), .B2(new_n934), .C1(new_n452), .C2(new_n762), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT46), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n776), .A2(G116), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n938), .B1(new_n936), .B2(new_n937), .C1(new_n939), .C2(new_n747), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G294), .A2(new_n774), .B1(new_n778), .B2(G97), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n220), .B2(new_n768), .C1(new_n758), .C2(new_n814), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n933), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n809), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n925), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n918), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n725), .A2(new_n208), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT88), .B1(new_n669), .B2(new_n671), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n673), .B(new_n670), .C1(new_n666), .C2(new_n668), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n680), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n678), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n615), .B(new_n621), .C1(new_n616), .C2(new_n655), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n626), .A2(new_n654), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT103), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT103), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n953), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n953), .A2(new_n964), .A3(new_n954), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT44), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n681), .B2(new_n961), .ZN(new_n971));
  INV_X1    g0771(.A(new_n961), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n679), .B1(new_n674), .B2(new_n675), .ZN(new_n973));
  OAI211_X1 g0773(.A(KEYINPUT44), .B(new_n972), .C1(new_n973), .C2(new_n678), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n677), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n663), .A2(G330), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n676), .A2(new_n680), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n979), .A2(new_n980), .A3(new_n973), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n979), .B1(new_n980), .B2(new_n973), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n719), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n966), .A2(new_n967), .B1(new_n971), .B2(new_n974), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(new_n677), .A3(new_n969), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n978), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n720), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n684), .B(KEYINPUT41), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n950), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n972), .B2(new_n953), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n973), .A2(KEYINPUT42), .A3(new_n961), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n565), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n961), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n615), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n655), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT104), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT43), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT43), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n993), .A2(new_n994), .B1(new_n998), .B2(new_n655), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT104), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n916), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n917), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n677), .A2(new_n972), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n916), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n948), .B1(new_n991), .B2(new_n1016), .ZN(G387));
  INV_X1    g0817(.A(new_n984), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n983), .A2(new_n719), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n684), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n686), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n739), .A2(new_n1021), .B1(new_n220), .B2(new_n683), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT110), .Z(new_n1023));
  NAND2_X1  g0823(.A1(new_n308), .A2(new_n201), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n686), .B(new_n273), .C1(new_n203), .C2(new_n218), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n737), .B1(new_n1025), .B2(new_n1026), .C1(new_n242), .C2(new_n273), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n727), .B1(new_n1028), .B2(new_n919), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n308), .A2(new_n774), .B1(new_n776), .B2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n779), .A2(new_n577), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n463), .C2(new_n766), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n812), .A2(G50), .B1(new_n783), .B2(G68), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n324), .C1(new_n747), .C2(new_n264), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G159), .C2(new_n786), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n321), .B1(new_n766), .B2(new_n456), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n812), .A2(G317), .B1(new_n783), .B2(G303), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n814), .B2(new_n764), .C1(new_n758), .C2(new_n781), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT48), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n776), .A2(G294), .B1(new_n779), .B2(G283), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1036), .B(new_n1045), .C1(G326), .C2(new_n748), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1035), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1029), .B1(new_n676), .B2(new_n790), .C1(new_n1048), .C2(new_n809), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1020), .B(new_n1049), .C1(new_n983), .C2(new_n949), .ZN(G393));
  OAI221_X1 g0850(.A(new_n919), .B1(new_n463), .B2(new_n234), .C1(new_n920), .C2(new_n253), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n726), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n758), .A2(new_n264), .B1(new_n330), .B2(new_n762), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n768), .A2(new_n218), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n203), .A2(new_n770), .B1(new_n766), .B2(new_n214), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G50), .C2(new_n774), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n324), .B1(new_n262), .B2(new_n761), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n748), .B2(G143), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n758), .A2(new_n939), .B1(new_n814), .B2(new_n762), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n339), .B1(new_n761), .B2(new_n527), .C1(new_n220), .C2(new_n766), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G303), .A2(new_n774), .B1(new_n776), .B2(G283), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n456), .B2(new_n768), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G322), .C2(new_n748), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1052), .B1(new_n1068), .B2(new_n734), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n961), .B2(new_n790), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n987), .A2(new_n684), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n984), .B1(new_n978), .B2(new_n986), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n976), .A2(new_n977), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n677), .B1(new_n985), .B2(new_n969), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n978), .A2(KEYINPUT111), .A3(new_n986), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1077), .A2(new_n950), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(KEYINPUT112), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1072), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n684), .A3(new_n987), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT112), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1077), .A2(new_n950), .A3(new_n1078), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1070), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1085), .ZN(G390));
  NAND4_X1  g0886(.A1(new_n717), .A2(new_n881), .A3(G330), .A4(new_n798), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n801), .A2(new_n883), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n881), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n863), .A2(new_n871), .B1(new_n1090), .B2(new_n865), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n900), .A2(new_n865), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n797), .A2(new_n432), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n655), .B(new_n1093), .C1(new_n696), .C2(new_n698), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n882), .B1(new_n1094), .B2(new_n883), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n843), .A2(new_n850), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n868), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n870), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n862), .A2(new_n895), .A3(new_n840), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n866), .B2(new_n884), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1087), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n718), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n439), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n887), .A2(new_n647), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n882), .B1(new_n718), .B2(new_n799), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n1087), .B1(new_n883), .B2(new_n801), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1094), .A2(new_n883), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1109), .A2(new_n1087), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n684), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1097), .A2(new_n1104), .A3(new_n950), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n731), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n726), .B1(new_n308), .B2(new_n806), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n764), .A2(new_n220), .B1(new_n761), .B2(new_n463), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n786), .B2(G283), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT113), .Z(new_n1124));
  OAI21_X1  g0924(.A(new_n339), .B1(new_n770), .B2(new_n214), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT114), .Z(new_n1126));
  AOI211_X1 g0926(.A(new_n1055), .B(new_n822), .C1(G116), .C2(new_n812), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n527), .C2(new_n747), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n289), .B1(new_n761), .B2(new_n1129), .C1(new_n824), .C2(new_n762), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n770), .A2(new_n264), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(KEYINPUT53), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G125), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1133), .B1(KEYINPUT53), .B2(new_n1132), .C1(new_n1134), .C2(new_n747), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n778), .A2(G50), .B1(new_n779), .B2(G159), .ZN(new_n1136));
  INV_X1    g0936(.A(G137), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n764), .C1(new_n758), .C2(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1124), .A2(new_n1128), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1121), .B1(new_n1140), .B2(new_n734), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1120), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1118), .A2(new_n1119), .A3(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(new_n1108), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1117), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT115), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n851), .A2(new_n862), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n1148));
  OAI21_X1  g0948(.A(G330), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT40), .B1(new_n875), .B2(new_n894), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n898), .A2(new_n904), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n270), .A2(new_n873), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n306), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n305), .A2(new_n270), .A3(new_n873), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1151), .A2(new_n1152), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(KEYINPUT115), .A3(new_n1159), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1163), .A3(new_n886), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n886), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1166));
  OAI211_X1 g0966(.A(KEYINPUT57), .B(new_n1145), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n684), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n886), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT116), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n872), .A2(new_n1172), .A3(new_n885), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n872), .B2(new_n885), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1163), .A3(new_n1161), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1145), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1168), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n778), .A2(G58), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n218), .B2(new_n770), .C1(new_n463), .C2(new_n764), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n321), .A2(new_n272), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n762), .A2(new_n220), .B1(new_n761), .B2(new_n426), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G68), .C2(new_n779), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n934), .B2(new_n747), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1181), .B(new_n1185), .C1(G116), .C2(new_n786), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT58), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT58), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1182), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n762), .A2(new_n1138), .B1(new_n761), .B2(new_n1137), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G132), .B2(new_n774), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1129), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n776), .A2(new_n1193), .B1(new_n779), .B2(G150), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(new_n1134), .C2(new_n758), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n748), .A2(G124), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n265), .B(new_n272), .C1(new_n766), .C2(new_n330), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n734), .B1(new_n1190), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1201), .B(new_n726), .C1(G50), .C2(new_n806), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1159), .B2(new_n731), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1177), .B2(new_n950), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1179), .A2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1115), .A2(new_n990), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n324), .B1(new_n264), .B2(new_n761), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1180), .B1(new_n201), .B2(new_n768), .C1(new_n330), .C2(new_n770), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(G128), .C2(new_n748), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT118), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n774), .A2(new_n1193), .B1(new_n812), .B2(G137), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n758), .B2(new_n824), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1031), .B1(new_n934), .B2(new_n762), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT117), .Z(new_n1215));
  OAI21_X1  g1015(.A(new_n339), .B1(new_n761), .B2(new_n220), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n764), .A2(new_n456), .B1(new_n770), .B2(new_n463), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G77), .C2(new_n778), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n527), .B2(new_n758), .C1(new_n452), .C2(new_n747), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1211), .A2(new_n1213), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n734), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n727), .B1(new_n203), .B2(new_n805), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n881), .C2(new_n732), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1113), .B2(new_n949), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1207), .A2(new_n1225), .ZN(G381));
  INV_X1    g1026(.A(G387), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(G384), .A2(G393), .A3(G381), .A4(G396), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OR3_X1    g1029(.A1(new_n1229), .A2(KEYINPUT119), .A3(G390), .ZN(new_n1230));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  INV_X1    g1031(.A(G375), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT119), .B1(new_n1229), .B2(G390), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(G407));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n653), .A3(new_n1231), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G390), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1080), .A2(KEYINPUT123), .A3(new_n1085), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(G387), .A3(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n794), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G387), .B1(new_n1085), .B2(new_n1080), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(KEYINPUT124), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G390), .A2(new_n1227), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1240), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G390), .A2(new_n1227), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1248), .B2(new_n1242), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n989), .B1(new_n1117), .B2(new_n1144), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1175), .A2(new_n1163), .A3(new_n1161), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n1166), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT120), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1171), .A2(new_n1164), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1203), .B1(new_n1256), .B2(new_n950), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1177), .A2(new_n1258), .A3(new_n1252), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1231), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G378), .B(new_n1204), .C1(new_n1168), .C2(new_n1178), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT121), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1108), .A2(new_n1113), .A3(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n684), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1115), .A2(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1206), .ZN(new_n1268));
  OR3_X1    g1068(.A1(G384), .A2(new_n1268), .A3(new_n1224), .ZN(new_n1269));
  OAI21_X1  g1069(.A(G384), .B1(new_n1224), .B2(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT121), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1261), .A2(new_n1262), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n653), .A2(G213), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1264), .A2(new_n1271), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1263), .A2(new_n1274), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1271), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(new_n1276), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1275), .A2(new_n1276), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1282), .B(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1271), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1281), .B1(new_n1277), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1251), .B1(new_n1280), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1275), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1263), .A2(new_n1274), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT125), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1263), .A2(new_n1297), .A3(new_n1294), .A4(new_n1274), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1272), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1285), .B(new_n1287), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1299), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1290), .B1(new_n1305), .B2(new_n1306), .ZN(G405));
  XNOR2_X1  g1107(.A(G375), .B(new_n1231), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1250), .A2(KEYINPUT127), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1250), .B1(KEYINPUT127), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1308), .A2(KEYINPUT127), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(new_n1278), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  OAI22_X1  g1114(.A1(new_n1309), .A2(new_n1310), .B1(new_n1278), .B2(new_n1312), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(G402));
endmodule


