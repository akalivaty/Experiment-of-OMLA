//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  AND2_X1   g000(.A1(KEYINPUT64), .A2(G146), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT64), .A2(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(G143), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT0), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n189), .A2(KEYINPUT65), .A3(new_n192), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n188), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n190), .A2(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n193), .A2(new_n194), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n205), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n211), .B1(new_n214), .B2(new_n194), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n191), .B1(new_n213), .B2(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT68), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n189), .A2(KEYINPUT68), .A3(new_n192), .A4(new_n217), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n210), .B1(G125), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT81), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(G224), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(G224), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n229), .A3(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT74), .ZN(new_n236));
  INV_X1    g050(.A(G107), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G104), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(G104), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n242), .A3(new_n237), .A4(G104), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(KEYINPUT4), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G101), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n239), .A2(new_n248), .A3(new_n241), .A4(new_n243), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(new_n245), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n244), .A2(new_n250), .A3(G101), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n245), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT76), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n235), .B(new_n247), .C1(new_n256), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n261));
  INV_X1    g075(.A(G119), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G116), .ZN(new_n263));
  INV_X1    g077(.A(new_n232), .ZN(new_n264));
  OAI211_X1 g078(.A(G113), .B(new_n263), .C1(new_n264), .C2(new_n261), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n264), .B2(new_n233), .ZN(new_n266));
  INV_X1    g080(.A(G104), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G107), .ZN(new_n268));
  OAI21_X1  g082(.A(G101), .B1(new_n240), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n249), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(G110), .B(G122), .Z(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n274), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n260), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(KEYINPUT6), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n253), .B1(new_n252), .B2(new_n255), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n257), .A2(KEYINPUT76), .A3(new_n258), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n246), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n271), .B1(new_n281), .B2(new_n235), .ZN(new_n282));
  NOR4_X1   g096(.A1(new_n282), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n276), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n276), .B1(new_n260), .B2(new_n272), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n231), .B(new_n278), .C1(new_n283), .C2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n223), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n225), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n290), .A2(KEYINPUT7), .B1(new_n227), .B2(G224), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n290), .B2(KEYINPUT7), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n222), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n274), .B(KEYINPUT8), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n266), .A2(new_n270), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n272), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n282), .B2(new_n276), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n288), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G210), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n288), .A2(new_n301), .A3(new_n299), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(KEYINPUT83), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n307), .A3(new_n302), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n194), .A2(G119), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT72), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n262), .B2(G128), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT24), .B(G110), .ZN(new_n313));
  INV_X1    g127(.A(G110), .ZN(new_n314));
  OR3_X1    g128(.A1(new_n262), .A2(KEYINPUT23), .A3(G128), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(new_n262), .B2(G128), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(G125), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(G146), .B(new_n321), .C1(new_n323), .C2(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n213), .A2(new_n322), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n323), .B2(new_n319), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n190), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n324), .ZN(new_n330));
  OAI221_X1 g144(.A(new_n330), .B1(new_n314), .B2(new_n317), .C1(new_n312), .C2(new_n313), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT22), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(G137), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G902), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n327), .A2(new_n331), .A3(new_n335), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT25), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(G234), .B2(new_n338), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n337), .A2(new_n344), .A3(new_n338), .A4(new_n339), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n337), .A2(new_n339), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n343), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G134), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n351), .B2(G137), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n353), .B(G131), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT66), .B1(new_n351), .B2(G137), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT11), .ZN(new_n358));
  INV_X1    g172(.A(new_n352), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT11), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT66), .B(new_n361), .C1(new_n351), .C2(G137), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n221), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n198), .A2(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n234), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n370), .A2(new_n200), .A3(new_n208), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n189), .A2(new_n192), .A3(new_n217), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT68), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n219), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n364), .B1(new_n378), .B2(new_n215), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT30), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n366), .A2(new_n381), .A3(new_n371), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n373), .B1(new_n383), .B2(new_n235), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G210), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n385), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT26), .B(G101), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT70), .B1(new_n384), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n235), .B1(new_n374), .B2(new_n379), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n372), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n372), .A2(new_n393), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n391), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n234), .B1(new_n380), .B2(new_n382), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n400), .B(new_n390), .C1(new_n401), .C2(new_n373), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n392), .A2(new_n398), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT71), .B1(new_n398), .B2(new_n399), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n397), .A2(new_n405), .A3(KEYINPUT29), .A4(new_n391), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n338), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G472), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n390), .B1(new_n395), .B2(new_n396), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n374), .A2(new_n379), .A3(KEYINPUT30), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n381), .B1(new_n366), .B2(new_n371), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n235), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n372), .A3(new_n391), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT31), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G472), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n384), .A2(KEYINPUT31), .A3(new_n391), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n338), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT32), .ZN(new_n419));
  INV_X1    g233(.A(new_n413), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n420), .B2(KEYINPUT31), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n415), .A4(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n350), .B1(new_n408), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G221), .B1(new_n427), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n367), .B(new_n247), .C1(new_n256), .C2(new_n259), .ZN(new_n430));
  INV_X1    g244(.A(new_n370), .ZN(new_n431));
  INV_X1    g245(.A(new_n216), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G128), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n378), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n270), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n437), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n430), .A2(new_n431), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(G110), .B(G140), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT73), .ZN(new_n444));
  INV_X1    g258(.A(G227), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n444), .B(new_n446), .Z(new_n447));
  AND2_X1   g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n430), .A2(new_n440), .A3(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n370), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n370), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n378), .A2(new_n215), .A3(new_n270), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT12), .B(new_n452), .C1(new_n438), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n377), .A2(new_n219), .B1(new_n432), .B2(new_n434), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n270), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n442), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n447), .B1(new_n461), .B2(KEYINPUT78), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n442), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  AOI221_X4 g278(.A(KEYINPUT79), .B1(new_n448), .B2(new_n450), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(KEYINPUT78), .ZN(new_n467));
  INV_X1    g281(.A(new_n447), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n448), .A2(new_n450), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G469), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G469), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n447), .B1(new_n450), .B2(new_n442), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n442), .A2(new_n460), .A3(new_n447), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n338), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n473), .B2(new_n338), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n429), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n323), .A2(G146), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n325), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n484), .A3(new_n325), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n386), .B2(G214), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n386), .A2(G143), .A3(G214), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT18), .A2(G131), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(G131), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n488), .A2(new_n360), .A3(new_n489), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(KEYINPUT17), .A3(G131), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n329), .A4(new_n324), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n267), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT85), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n496), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT19), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n322), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n213), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n324), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n501), .B1(new_n493), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n480), .B(new_n338), .C1(new_n503), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n493), .A2(new_n509), .ZN(new_n514));
  INV_X1    g328(.A(new_n501), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n493), .A2(new_n499), .A3(new_n502), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(KEYINPUT86), .A3(new_n480), .A4(new_n338), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n519), .A3(KEYINPUT20), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n501), .B1(new_n493), .B2(new_n499), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n338), .B1(new_n503), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G475), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n512), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n202), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n194), .A2(G143), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G134), .ZN(new_n530));
  XNOR2_X1  g344(.A(G128), .B(G143), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n351), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n530), .B2(new_n532), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G122), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G116), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(G116), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n237), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n539), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT89), .B1(new_n539), .B2(KEYINPUT14), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT88), .B(new_n540), .C1(new_n538), .C2(new_n544), .ZN(new_n549));
  AND4_X1   g363(.A1(new_n543), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n536), .B(new_n542), .C1(new_n550), .C2(new_n237), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n541), .B(new_n237), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n531), .A2(KEYINPUT13), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(G134), .C1(KEYINPUT13), .C2(new_n527), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n554), .A3(new_n532), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n427), .A2(new_n342), .A3(G953), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n555), .A3(new_n557), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n338), .ZN(new_n562));
  INV_X1    g376(.A(G478), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n562), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(G234), .A2(G237), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(G952), .A3(new_n227), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT21), .B(G898), .Z(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(G902), .A3(G953), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n526), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n309), .A2(new_n425), .A3(new_n479), .A4(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  NAND4_X1  g388(.A1(new_n288), .A2(KEYINPUT90), .A3(new_n301), .A4(new_n299), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n306), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT90), .B1(new_n300), .B2(new_n302), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n304), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n559), .A2(new_n580), .A3(new_n560), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n559), .B2(new_n560), .ZN(new_n582));
  OAI211_X1 g396(.A(G478), .B(new_n338), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT91), .B(G478), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n562), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n526), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n579), .A2(new_n571), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n421), .A2(new_n415), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G472), .ZN(new_n590));
  INV_X1    g404(.A(new_n350), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n418), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n429), .B(new_n592), .C1(new_n472), .C2(new_n478), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT92), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n594), .B(new_n596), .ZN(G6));
  INV_X1    g411(.A(new_n526), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n565), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n579), .A2(new_n571), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n593), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G107), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NOR2_X1   g417(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n332), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n348), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n346), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n590), .A2(new_n418), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n309), .A2(new_n479), .A3(new_n572), .A4(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT37), .B(G110), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  XOR2_X1   g426(.A(new_n567), .B(KEYINPUT93), .Z(new_n613));
  INV_X1    g427(.A(G900), .ZN(new_n614));
  INV_X1    g428(.A(new_n569), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n599), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n607), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n408), .B2(new_n424), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n479), .A2(new_n578), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n576), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT90), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n303), .A2(new_n624), .A3(new_n304), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n626), .A2(KEYINPUT94), .A3(new_n479), .A4(new_n617), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G128), .ZN(G30));
  NAND2_X1  g443(.A1(new_n305), .A2(new_n308), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n424), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n391), .B1(new_n401), .B2(new_n373), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n394), .A2(new_n372), .A3(new_n390), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n338), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n416), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n306), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n526), .A2(new_n565), .ZN(new_n640));
  NOR4_X1   g454(.A1(new_n638), .A2(new_n639), .A3(new_n607), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n616), .B(KEYINPUT39), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n479), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT40), .Z(new_n648));
  NAND3_X1  g462(.A1(new_n632), .A2(KEYINPUT95), .A3(new_n641), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n644), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT96), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n644), .A2(new_n648), .A3(new_n652), .A4(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n202), .ZN(G45));
  INV_X1    g469(.A(new_n616), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n526), .A2(new_n586), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT97), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n526), .A2(new_n586), .A3(new_n659), .A4(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n479), .A2(new_n578), .A3(new_n619), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n338), .B1(new_n474), .B2(new_n475), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G469), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n476), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n665), .B1(new_n668), .B2(new_n429), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n667), .A2(KEYINPUT98), .A3(new_n428), .A4(new_n476), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n425), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n588), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NAND2_X1  g490(.A1(new_n600), .A2(new_n673), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  INV_X1    g492(.A(new_n671), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n626), .A3(new_n572), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NOR2_X1   g495(.A1(new_n671), .A2(new_n592), .ZN(new_n682));
  INV_X1    g496(.A(new_n640), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n570), .A3(new_n578), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  NOR2_X1   g499(.A1(new_n661), .A2(new_n608), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n578), .A3(new_n669), .A4(new_n670), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G125), .ZN(G27));
  AOI21_X1  g502(.A(new_n639), .B1(new_n305), .B2(new_n308), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n469), .A2(G469), .A3(new_n470), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n473), .A2(new_n338), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT99), .Z(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n476), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n428), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n425), .A3(new_n662), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT42), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n360), .ZN(G33));
  NAND4_X1  g511(.A1(new_n689), .A2(new_n425), .A3(new_n617), .A4(new_n694), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n351), .ZN(G36));
  AND2_X1   g517(.A1(new_n590), .A2(new_n418), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n618), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT103), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT102), .B1(new_n598), .B2(new_n586), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT43), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n706), .A2(KEYINPUT44), .A3(new_n708), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(new_n689), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n476), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n469), .A2(KEYINPUT45), .A3(new_n470), .ZN(new_n715));
  INV_X1    g529(.A(new_n464), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n463), .B1(new_n442), .B2(new_n460), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n447), .ZN(new_n718));
  INV_X1    g532(.A(new_n470), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT79), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n469), .A2(new_n466), .A3(new_n470), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(G469), .B(new_n715), .C1(new_n722), .C2(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n692), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n714), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n692), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n429), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n646), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(KEYINPUT101), .A3(new_n646), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n713), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G137), .ZN(G39));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT105), .B1(new_n728), .B2(new_n735), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n735), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n728), .A2(new_n735), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n728), .A2(KEYINPUT104), .A3(new_n735), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n736), .A2(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n408), .A2(new_n424), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n591), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n662), .A3(new_n689), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G140), .ZN(G42));
  AND2_X1   g560(.A1(new_n708), .A2(new_n613), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n630), .B(KEYINPUT38), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n639), .A4(new_n682), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n679), .A2(new_n689), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n747), .A3(new_n609), .ZN(new_n754));
  INV_X1    g568(.A(new_n638), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n752), .A2(new_n350), .A3(new_n567), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n598), .A3(new_n585), .A4(new_n583), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n751), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT115), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n751), .A2(new_n760), .A3(new_n757), .A4(new_n754), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n592), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n747), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n668), .A2(new_n428), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n689), .B(new_n764), .C1(new_n742), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n766), .A3(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n227), .A2(G952), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n753), .A2(new_n747), .A3(new_n425), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT48), .Z(new_n770));
  INV_X1    g584(.A(new_n587), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n768), .B(new_n770), .C1(new_n771), .C2(new_n756), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n758), .B(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT51), .B1(new_n775), .B2(new_n766), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n663), .A2(new_n687), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n622), .B2(new_n627), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n579), .A2(new_n640), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n607), .A2(new_n616), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT112), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n755), .A3(new_n694), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n780), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n781), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n780), .A2(new_n628), .A3(new_n788), .A4(new_n786), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n779), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n628), .A2(new_n788), .A3(new_n786), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n782), .A2(new_n780), .A3(new_n786), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n662), .A2(new_n694), .A3(new_n704), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n473), .B1(new_n720), .B2(new_n721), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n743), .B(new_n428), .C1(new_n797), .C2(new_n477), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n526), .A2(new_n565), .A3(new_n616), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n607), .A3(new_n689), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n700), .B2(new_n701), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n674), .A2(new_n677), .A3(new_n680), .A4(new_n684), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n696), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n801), .B(KEYINPUT110), .C1(new_n700), .C2(new_n701), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(new_n599), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n309), .A2(new_n810), .A3(new_n570), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n305), .A2(new_n306), .A3(new_n308), .A4(new_n570), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT108), .B1(new_n813), .B2(new_n599), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n593), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n610), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n763), .B(new_n428), .C1(new_n797), .C2(new_n477), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n813), .A3(new_n587), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n428), .B(new_n572), .C1(new_n797), .C2(new_n477), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n672), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n593), .A2(new_n309), .A3(new_n570), .A4(new_n771), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT107), .A3(new_n573), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT109), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n816), .A2(new_n826), .A3(KEYINPUT109), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n809), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(KEYINPUT111), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n805), .B1(new_n802), .B2(new_n803), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n807), .A2(new_n808), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n816), .A2(new_n826), .A3(KEYINPUT109), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n827), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n778), .B(new_n795), .C1(new_n831), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n792), .A2(new_n793), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n764), .A2(new_n578), .A3(new_n679), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n790), .A2(KEYINPUT53), .A3(new_n794), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n830), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n778), .B1(new_n835), .B2(new_n839), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n777), .A2(new_n841), .A3(new_n842), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(G952), .B2(G953), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n598), .A2(new_n586), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n851), .A2(new_n350), .A3(new_n639), .A4(new_n429), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT106), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n755), .B1(new_n853), .B2(KEYINPUT49), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n668), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n748), .A2(new_n852), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n850), .A2(new_n857), .ZN(G75));
  OAI21_X1  g672(.A(new_n278), .B1(new_n283), .B2(new_n287), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(new_n231), .Z(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT55), .ZN(new_n861));
  INV_X1    g675(.A(G210), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n862), .B(new_n338), .C1(new_n844), .C2(new_n846), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n863), .B2(KEYINPUT56), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n227), .A2(G952), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n844), .A2(new_n846), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(G210), .A3(G902), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  INV_X1    g683(.A(new_n861), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n864), .A2(new_n874), .A3(new_n871), .A4(new_n866), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(G51));
  XOR2_X1   g690(.A(new_n692), .B(KEYINPUT57), .Z(new_n877));
  AOI21_X1  g691(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n847), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n474), .A2(new_n475), .ZN(new_n882));
  OAI211_X1 g696(.A(KEYINPUT117), .B(new_n877), .C1(new_n847), .C2(new_n878), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n867), .A2(G902), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(new_n723), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n865), .B1(new_n884), .B2(new_n886), .ZN(G54));
  NAND4_X1  g701(.A1(new_n867), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  INV_X1    g703(.A(new_n518), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n865), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G60));
  NOR2_X1   g708(.A1(new_n581), .A2(new_n582), .ZN(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n563), .A2(new_n338), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n847), .B2(new_n878), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n841), .B2(new_n848), .ZN(new_n901));
  INV_X1    g715(.A(new_n895), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n866), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT60), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n867), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n347), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n867), .A2(new_n605), .A3(new_n906), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n866), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G66));
  NAND2_X1  g727(.A1(new_n568), .A2(G224), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(G953), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n805), .B1(new_n828), .B2(new_n829), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(G953), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT120), .Z(new_n918));
  OAI21_X1  g732(.A(new_n859), .B1(G898), .B2(new_n227), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  INV_X1    g734(.A(new_n647), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n599), .A2(new_n587), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n425), .A3(new_n689), .A4(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n733), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n651), .A2(new_n653), .A3(new_n782), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT62), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n925), .B2(KEYINPUT62), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n745), .B(new_n924), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n651), .A2(new_n931), .A3(new_n653), .A4(new_n782), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n227), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n505), .A2(new_n507), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT121), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n383), .B(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n445), .B2(new_n614), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n579), .A2(new_n672), .A3(new_n640), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n732), .B(new_n731), .C1(new_n713), .C2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n702), .A2(new_n696), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n745), .A2(new_n949), .A3(new_n227), .A4(new_n782), .ZN(new_n950));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n951), .A3(new_n939), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n941), .A2(new_n944), .A3(new_n945), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n927), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(new_n934), .A3(new_n745), .A4(new_n924), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n939), .B1(new_n957), .B2(new_n227), .ZN(new_n958));
  INV_X1    g772(.A(new_n952), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n943), .B(new_n942), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n953), .A2(new_n960), .ZN(G72));
  INV_X1    g775(.A(new_n916), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT126), .Z(new_n967));
  AOI21_X1  g781(.A(new_n634), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n392), .A2(new_n402), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n413), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n838), .A2(new_n840), .A3(new_n966), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n745), .A2(new_n949), .A3(new_n782), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n974), .B2(new_n962), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n384), .A3(new_n390), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n976), .A3(new_n866), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n968), .A2(new_n977), .ZN(G57));
endmodule


