//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1046, new_n1047;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT94), .ZN(new_n203));
  XOR2_X1   g002(.A(G169gat), .B(G197gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT12), .ZN(new_n208));
  INV_X1    g007(.A(new_n206), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n205), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT12), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G229gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(KEYINPUT14), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT15), .A4(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT15), .B1(new_n219), .B2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT14), .ZN(new_n226));
  NAND2_X1  g025(.A1(G29gat), .A2(G36gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n221), .A3(KEYINPUT15), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n215), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n222), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(G1gat), .ZN(new_n235));
  OAI21_X1  g034(.A(G8gat), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n233), .ZN(new_n237));
  INV_X1    g036(.A(G8gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n237), .B(new_n238), .C1(G1gat), .C2(new_n231), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT96), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT96), .B1(new_n236), .B2(new_n239), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n230), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n221), .A3(new_n227), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n228), .A3(new_n215), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n222), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n236), .A2(new_n239), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n245), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI211_X1 g054(.A(KEYINPUT95), .B(new_n240), .C1(new_n246), .C2(new_n252), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n214), .B(new_n244), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT97), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n213), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n252), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n251), .B1(new_n250), .B2(new_n222), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT95), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n253), .A2(new_n245), .A3(new_n254), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT18), .A3(new_n214), .A4(new_n244), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n254), .A2(KEYINPUT96), .ZN(new_n269));
  INV_X1    g068(.A(new_n243), .ZN(new_n270));
  INV_X1    g069(.A(new_n230), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n244), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n214), .B(KEYINPUT13), .Z(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n268), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n257), .A2(new_n258), .B1(new_n273), .B2(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT97), .B1(new_n257), .B2(new_n258), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n278), .B(new_n268), .C1(new_n279), .C2(new_n213), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT36), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT26), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT28), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n292), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n302), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n311), .B(new_n312), .C1(new_n313), .C2(KEYINPUT64), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n295), .A2(KEYINPUT64), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n308), .B(new_n309), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(new_n307), .B2(new_n292), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n287), .A2(KEYINPUT23), .A3(new_n289), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n315), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n311), .A3(new_n312), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT66), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(new_n320), .A3(new_n322), .A4(new_n325), .ZN(new_n326));
  AOI221_X4 g125(.A(KEYINPUT67), .B1(new_n317), .B2(new_n318), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n317), .A2(new_n318), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n306), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G134gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342));
  NAND2_X1  g141(.A1(G113gat), .A2(G120gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n333), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n338), .A2(new_n344), .A3(KEYINPUT70), .A4(new_n345), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n336), .A3(new_n342), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(new_n343), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n348), .A2(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G227gat), .ZN(new_n358));
  INV_X1    g157(.A(G233gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n348), .A2(new_n349), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n306), .B(new_n363), .C1(new_n327), .C2(new_n331), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n360), .A4(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT73), .B(KEYINPUT33), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT74), .ZN(new_n374));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n364), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n358), .B2(new_n359), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n379), .B(KEYINPUT34), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  INV_X1    g180(.A(new_n371), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AND4_X1   g182(.A1(new_n381), .A2(new_n369), .A3(KEYINPUT32), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT32), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n367), .B2(new_n368), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n381), .B1(new_n386), .B2(new_n383), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n377), .B(new_n380), .C1(new_n384), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT75), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n381), .A3(new_n383), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n380), .B1(new_n393), .B2(new_n377), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n283), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n377), .B1(new_n384), .B2(new_n387), .ZN(new_n396));
  INV_X1    g195(.A(new_n380), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(KEYINPUT36), .A3(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G1gat), .B(G29gat), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G141gat), .ZN(new_n406));
  INV_X1    g205(.A(G148gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409));
  AND2_X1   g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT2), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n415), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G155gat), .ZN(new_n418));
  INV_X1    g217(.A(G162gat), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT2), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(G141gat), .A2(G148gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n410), .A2(new_n413), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n420), .B(new_n423), .C1(new_n424), .C2(new_n415), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n356), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n361), .A2(KEYINPUT83), .A3(new_n362), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n361), .B2(new_n362), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n426), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT5), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n425), .A3(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT4), .B1(new_n439), .B2(new_n363), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n356), .A2(new_n441), .A3(new_n426), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n363), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n356), .A2(KEYINPUT83), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n425), .A3(KEYINPUT3), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n417), .B2(new_n425), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n448), .B2(new_n447), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n446), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(new_n434), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n443), .A2(new_n452), .A3(KEYINPUT85), .A4(new_n434), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n435), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n438), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT84), .B1(new_n417), .B2(new_n425), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n441), .A3(new_n356), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n428), .B2(new_n441), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n434), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT6), .B(new_n405), .C1(new_n457), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n455), .A2(new_n456), .ZN(new_n468));
  INV_X1    g267(.A(new_n435), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n466), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n404), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n405), .B1(new_n457), .B2(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n467), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n306), .B(new_n479), .C1(new_n327), .C2(new_n331), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n304), .B1(new_n297), .B2(new_n299), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n324), .A2(new_n326), .B1(new_n318), .B2(new_n317), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n478), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(G211gat), .A2(G218gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G211gat), .A2(G218gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT76), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT76), .ZN(new_n490));
  INV_X1    g289(.A(new_n488), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n486), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(G197gat), .A2(G204gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT22), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n493), .A2(KEYINPUT77), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n494), .A2(new_n495), .B1(new_n497), .B2(new_n488), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n492), .B(new_n489), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT78), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT78), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n485), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n482), .A2(new_n483), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n479), .ZN(new_n510));
  INV_X1    g309(.A(new_n331), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n483), .A2(new_n328), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n482), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n479), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n510), .B(new_n506), .C1(new_n513), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G8gat), .B(G36gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G64gat), .B(G92gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  NAND3_X1  g320(.A1(new_n508), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n522), .A2(KEYINPUT30), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n518), .ZN(new_n525));
  INV_X1    g324(.A(new_n521), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT80), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT80), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n528), .B(new_n521), .C1(new_n508), .C2(new_n518), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n523), .A2(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n477), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n515), .B1(new_n493), .B2(new_n499), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n501), .A2(new_n489), .A3(new_n492), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT3), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n460), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT3), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n439), .A3(KEYINPUT86), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n450), .A2(new_n515), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n500), .A2(new_n503), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT78), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n537), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G228gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G22gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n506), .A2(new_n553), .A3(new_n542), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n539), .B1(new_n543), .B2(KEYINPUT29), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n549), .B1(new_n555), .B2(new_n432), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n559));
  XNOR2_X1  g358(.A(G78gat), .B(G106gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G50gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n550), .A2(new_n557), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G22gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n558), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n559), .A2(new_n569), .A3(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n559), .B2(new_n562), .ZN(new_n572));
  INV_X1    g371(.A(new_n562), .ZN(new_n573));
  AOI211_X1 g372(.A(KEYINPUT89), .B(new_n573), .C1(new_n558), .C2(KEYINPUT88), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n567), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n532), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n467), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n457), .B2(new_n466), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT92), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n404), .B(KEYINPUT91), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT6), .B1(new_n585), .B2(new_n404), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n578), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n526), .B1(new_n525), .B2(KEYINPUT37), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n525), .A2(KEYINPUT37), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n510), .B1(new_n513), .B2(new_n517), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n593), .B2(new_n506), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n507), .B1(new_n480), .B2(new_n484), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n522), .B1(new_n596), .B2(new_n589), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n576), .B1(new_n587), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n530), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n433), .ZN(new_n602));
  INV_X1    g401(.A(new_n434), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n434), .B1(new_n462), .B2(new_n452), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n582), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT40), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n604), .A2(new_n606), .A3(new_n605), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n612), .A2(new_n613), .A3(new_n609), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n525), .A2(new_n526), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n528), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n525), .A2(KEYINPUT80), .A3(new_n526), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n522), .B(KEYINPUT30), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT90), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n601), .A2(new_n615), .A3(new_n621), .A4(new_n584), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n599), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n400), .A2(new_n577), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n586), .A2(new_n475), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n530), .B1(new_n625), .B2(new_n467), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n571), .A2(new_n575), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n398), .A2(new_n626), .A3(new_n627), .A4(new_n388), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n398), .A2(new_n627), .A3(new_n388), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n601), .A2(new_n621), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n584), .A2(new_n586), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n578), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n629), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n282), .B1(new_n624), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n477), .ZN(new_n637));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n418), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G71gat), .A2(G78gat), .ZN(new_n643));
  OR2_X1    g442(.A1(G71gat), .A2(G78gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT9), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(G57gat), .A2(G64gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(G57gat), .A2(G64gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(KEYINPUT99), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650));
  AND2_X1   g449(.A1(G57gat), .A2(G64gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(G57gat), .A2(G64gat), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n646), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n647), .A2(KEYINPUT9), .A3(new_n648), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n656));
  OR3_X1    g455(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .A4(new_n643), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT21), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n269), .A2(new_n270), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT21), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G231gat), .A2(G233gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G127gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n335), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n664), .A3(new_n665), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n642), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n672), .A2(new_n674), .A3(new_n642), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT7), .ZN(new_n679));
  OAI211_X1 g478(.A(G85gat), .B(G92gat), .C1(new_n679), .C2(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g479(.A1(G85gat), .A2(G92gat), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT7), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G99gat), .B(G106gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(G99gat), .A2(G106gat), .ZN(new_n686));
  INV_X1    g485(.A(G85gat), .ZN(new_n687));
  INV_X1    g486(.A(G92gat), .ZN(new_n688));
  AOI22_X1  g487(.A1(KEYINPUT8), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n685), .B1(new_n684), .B2(new_n689), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n230), .ZN(new_n694));
  NAND3_X1  g493(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  INV_X1    g495(.A(new_n693), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n253), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT103), .B(new_n693), .C1(new_n246), .C2(new_n252), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n694), .B(new_n695), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(G190gat), .B(G218gat), .Z(new_n701));
  OR2_X1    g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  XNOR2_X1  g502(.A(G134gat), .B(G162gat), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n704), .B(new_n705), .Z(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT104), .Z(new_n707));
  AND3_X1   g506(.A1(new_n702), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n702), .A2(new_n703), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n659), .B1(new_n691), .B2(new_n692), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n684), .A2(new_n689), .ZN(new_n713));
  INV_X1    g512(.A(new_n685), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n715), .A2(new_n658), .A3(new_n654), .A4(new_n690), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT10), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n693), .A2(new_n660), .A3(KEYINPUT10), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(G230gat), .A2(G233gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n712), .B2(new_n716), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(G120gat), .B(G148gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(G176gat), .B(G204gat), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n725), .B(new_n726), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n727), .ZN(new_n729));
  INV_X1    g528(.A(new_n721), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n718), .B2(new_n719), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n678), .A2(new_n711), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT106), .Z(new_n740));
  NAND3_X1  g539(.A1(new_n636), .A2(new_n637), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g541(.A1(new_n636), .A2(new_n740), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n631), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT16), .B(G8gat), .Z(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n238), .B2(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1325gat));
  OAI21_X1  g550(.A(G15gat), .B1(new_n743), .B2(new_n400), .ZN(new_n752));
  INV_X1    g551(.A(G15gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n398), .A2(new_n388), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n636), .A2(new_n753), .A3(new_n755), .A4(new_n740), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(G1326gat));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n743), .B2(new_n627), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n636), .A2(KEYINPUT107), .A3(new_n576), .A4(new_n740), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT43), .B(G22gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1327gat));
  NOR3_X1   g562(.A1(new_n678), .A2(new_n711), .A3(new_n737), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n636), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n224), .A3(new_n637), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT45), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n711), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n626), .A2(new_n627), .ZN(new_n770));
  AOI221_X4 g569(.A(new_n770), .B1(new_n599), .B2(new_n622), .C1(new_n395), .C2(new_n399), .ZN(new_n771));
  INV_X1    g570(.A(new_n634), .ZN(new_n772));
  INV_X1    g571(.A(new_n630), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(new_n773), .B1(new_n628), .B2(KEYINPUT35), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n769), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776));
  INV_X1    g575(.A(new_n677), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n675), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n676), .A2(KEYINPUT108), .A3(new_n677), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(new_n282), .A3(new_n737), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n577), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n532), .A2(KEYINPUT109), .A3(new_n576), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n400), .A2(new_n623), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n711), .B1(new_n786), .B2(new_n635), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n775), .B(new_n782), .C1(new_n787), .C2(KEYINPUT44), .ZN(new_n788));
  OAI21_X1  g587(.A(G29gat), .B1(new_n788), .B2(new_n477), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n767), .A2(new_n789), .ZN(G1328gat));
  INV_X1    g589(.A(new_n631), .ZN(new_n791));
  AOI21_X1  g590(.A(G36gat), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n765), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G36gat), .B1(new_n788), .B2(new_n631), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1329gat));
  OAI21_X1  g596(.A(G43gat), .B1(new_n788), .B2(new_n400), .ZN(new_n798));
  INV_X1    g597(.A(G43gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n765), .A2(new_n799), .A3(new_n755), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(KEYINPUT47), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1330gat));
  OAI21_X1  g604(.A(KEYINPUT111), .B1(new_n788), .B2(new_n627), .ZN(new_n806));
  INV_X1    g605(.A(new_n769), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n624), .B2(new_n635), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n398), .A2(KEYINPUT36), .A3(new_n388), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT36), .B1(new_n398), .B2(new_n388), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n623), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n784), .A2(new_n785), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n628), .A2(KEYINPUT35), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n634), .A2(new_n630), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n708), .A2(new_n710), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n808), .B1(new_n817), .B2(new_n768), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n576), .A4(new_n782), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n806), .A2(new_n820), .A3(G50gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT48), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n627), .A2(G50gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n765), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G50gat), .B1(new_n788), .B2(new_n627), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n765), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n822), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(G1331gat));
  INV_X1    g629(.A(new_n678), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n831), .A2(new_n816), .A3(new_n281), .A4(new_n738), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n815), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n637), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G57gat), .ZN(G1332gat));
  AND3_X1   g634(.A1(new_n815), .A2(new_n791), .A3(new_n832), .ZN(new_n836));
  NOR2_X1   g635(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n837));
  AND2_X1   g636(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n840), .B(new_n841), .ZN(G1333gat));
  NAND4_X1  g641(.A1(new_n833), .A2(G71gat), .A3(new_n399), .A4(new_n395), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n754), .B(KEYINPUT113), .Z(new_n844));
  AND2_X1   g643(.A1(new_n833), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n845), .B2(G71gat), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g646(.A1(new_n833), .A2(new_n576), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g648(.A1(new_n678), .A2(new_n281), .A3(new_n738), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n775), .B(new_n850), .C1(new_n787), .C2(KEYINPUT44), .ZN(new_n851));
  OAI21_X1  g650(.A(G85gat), .B1(new_n851), .B2(new_n477), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n678), .A2(new_n281), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n815), .A2(new_n816), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n787), .A2(KEYINPUT51), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n637), .A2(new_n687), .A3(new_n737), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n852), .B1(new_n859), .B2(new_n860), .ZN(G1336gat));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n851), .B2(new_n631), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n791), .A4(new_n850), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(G92gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n631), .A2(G92gat), .A3(new_n738), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G92gat), .B1(new_n851), .B2(new_n631), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n855), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT51), .B1(new_n787), .B2(new_n853), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(G1337gat));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n851), .B2(new_n400), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G99gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n400), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n754), .A2(G99gat), .A3(new_n738), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT116), .Z(new_n880));
  OAI22_X1  g679(.A1(new_n877), .A2(new_n878), .B1(new_n859), .B2(new_n880), .ZN(G1338gat));
  NOR3_X1   g680(.A1(new_n627), .A2(G106gat), .A3(new_n738), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n858), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G106gat), .B1(new_n851), .B2(new_n627), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1339gat));
  NAND3_X1  g688(.A1(new_n718), .A2(new_n719), .A3(new_n730), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n722), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n727), .B1(new_n731), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(KEYINPUT55), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n728), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT55), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT117), .B(KEYINPUT55), .C1(new_n891), .C2(new_n893), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n280), .B2(new_n277), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n259), .A2(new_n268), .A3(new_n213), .A4(new_n275), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n271), .B1(new_n269), .B2(new_n270), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n265), .B2(new_n266), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n905), .A2(new_n214), .B1(new_n273), .B2(new_n274), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n207), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n737), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n711), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n903), .A2(new_n907), .ZN(new_n910));
  INV_X1    g709(.A(new_n901), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n816), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n781), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n739), .A2(new_n281), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT118), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n281), .ZN(new_n916));
  INV_X1    g715(.A(new_n908), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n816), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n816), .A2(new_n910), .A3(new_n911), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n780), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n921));
  INV_X1    g720(.A(new_n914), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n915), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n631), .A2(new_n637), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n773), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n282), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(new_n339), .ZN(G1340gat));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n738), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(new_n340), .ZN(G1341gat));
  OAI21_X1  g730(.A(G127gat), .B1(new_n927), .B2(new_n780), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n678), .A2(new_n335), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n927), .B2(new_n933), .ZN(G1342gat));
  OR2_X1    g733(.A1(new_n927), .A2(new_n711), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G134gat), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT56), .B1(new_n935), .B2(G134gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(G134gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(KEYINPUT119), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT119), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n936), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(G1343gat));
  AOI21_X1  g741(.A(new_n925), .B1(new_n395), .B2(new_n399), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n915), .A2(new_n923), .A3(new_n576), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n897), .A2(new_n898), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n728), .A3(new_n894), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n277), .B2(new_n280), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n711), .B1(new_n951), .B2(new_n908), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT120), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n954), .B(new_n711), .C1(new_n951), .C2(new_n908), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(new_n912), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n831), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n948), .B1(new_n957), .B2(new_n922), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n944), .B1(new_n947), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n406), .B1(new_n960), .B2(new_n281), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n915), .A3(new_n576), .A4(new_n923), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n281), .A2(new_n406), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n961), .A2(KEYINPUT58), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(KEYINPUT121), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n967), .B1(new_n962), .B2(new_n963), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g768(.A(KEYINPUT122), .B(KEYINPUT58), .C1(new_n961), .C2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n958), .B1(new_n945), .B2(new_n946), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n972), .A2(new_n282), .A3(new_n944), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n968), .B(new_n966), .C1(new_n973), .C2(new_n406), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT122), .B1(new_n974), .B2(KEYINPUT58), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n965), .B1(new_n971), .B2(new_n975), .ZN(G1344gat));
  INV_X1    g775(.A(new_n962), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n407), .A3(new_n737), .ZN(new_n978));
  XOR2_X1   g777(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n979));
  AND2_X1   g778(.A1(new_n740), .A2(new_n282), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n678), .B1(new_n912), .B2(new_n952), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n576), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n946), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n924), .A2(KEYINPUT57), .A3(new_n576), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n985), .A2(new_n737), .A3(new_n943), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n979), .B1(new_n986), .B2(G148gat), .ZN(new_n987));
  AOI211_X1 g786(.A(KEYINPUT59), .B(new_n407), .C1(new_n960), .C2(new_n737), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n978), .B1(new_n987), .B2(new_n988), .ZN(G1345gat));
  NOR2_X1   g788(.A1(new_n962), .A2(new_n831), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  AOI21_X1  g790(.A(G155gat), .B1(new_n990), .B2(KEYINPUT124), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n780), .A2(new_n418), .ZN(new_n993));
  AOI22_X1  g792(.A1(new_n991), .A2(new_n992), .B1(new_n960), .B2(new_n993), .ZN(G1346gat));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n419), .A3(new_n816), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n972), .A2(new_n711), .A3(new_n944), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(new_n419), .ZN(G1347gat));
  NOR2_X1   g796(.A1(new_n631), .A2(new_n637), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n844), .A2(new_n627), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(new_n924), .ZN(new_n1000));
  OAI21_X1  g799(.A(G169gat), .B1(new_n1000), .B2(new_n282), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n924), .A2(new_n773), .A3(new_n998), .ZN(new_n1003));
  INV_X1    g802(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n282), .A2(G169gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR4_X1   g805(.A1(new_n1003), .A2(KEYINPUT125), .A3(G169gat), .A4(new_n282), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n1001), .B(new_n1010), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1348gat));
  OAI21_X1  g811(.A(G176gat), .B1(new_n1000), .B2(new_n738), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1004), .A2(new_n286), .A3(new_n737), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1349gat));
  OAI21_X1  g814(.A(G183gat), .B1(new_n1000), .B2(new_n780), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1004), .A2(new_n301), .A3(new_n678), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n302), .A3(new_n816), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n999), .A2(new_n816), .A3(new_n924), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1022));
  AND4_X1   g821(.A1(KEYINPUT127), .A2(new_n1021), .A3(new_n1022), .A4(G190gat), .ZN(new_n1023));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n302), .B1(new_n1024), .B2(KEYINPUT61), .ZN(new_n1025));
  AOI22_X1  g824(.A1(new_n1021), .A2(new_n1025), .B1(KEYINPUT127), .B2(new_n1022), .ZN(new_n1026));
  OAI21_X1  g825(.A(new_n1020), .B1(new_n1023), .B2(new_n1026), .ZN(G1351gat));
  NAND2_X1  g826(.A1(new_n400), .A2(new_n998), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n1029), .A2(new_n924), .A3(new_n576), .ZN(new_n1030));
  INV_X1    g829(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g830(.A(G197gat), .B1(new_n1031), .B2(new_n281), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1028), .B1(new_n983), .B2(new_n984), .ZN(new_n1033));
  AND2_X1   g832(.A1(new_n281), .A2(G197gat), .ZN(new_n1034));
  AOI21_X1  g833(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(G1352gat));
  NOR3_X1   g834(.A1(new_n1030), .A2(G204gat), .A3(new_n738), .ZN(new_n1036));
  XNOR2_X1  g835(.A(new_n1036), .B(KEYINPUT62), .ZN(new_n1037));
  INV_X1    g836(.A(new_n1033), .ZN(new_n1038));
  OAI21_X1  g837(.A(G204gat), .B1(new_n1038), .B2(new_n738), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1037), .A2(new_n1039), .ZN(G1353gat));
  OR3_X1    g839(.A1(new_n1030), .A2(G211gat), .A3(new_n831), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1033), .A2(new_n678), .ZN(new_n1042));
  AND3_X1   g841(.A1(new_n1042), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1043));
  AOI21_X1  g842(.A(KEYINPUT63), .B1(new_n1042), .B2(G211gat), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G1354gat));
  OAI21_X1  g844(.A(G218gat), .B1(new_n1038), .B2(new_n711), .ZN(new_n1046));
  OR3_X1    g845(.A1(new_n1030), .A2(G218gat), .A3(new_n711), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(G1355gat));
endmodule


