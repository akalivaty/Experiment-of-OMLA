//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT74), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n202), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT69), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(new_n219), .B2(KEYINPUT69), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(KEYINPUT69), .B(new_n222), .C1(new_n219), .C2(new_n220), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n217), .A2(new_n226), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT39), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n236));
  OAI211_X1 g035(.A(new_n235), .B(new_n226), .C1(new_n217), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n228), .A2(KEYINPUT4), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n217), .B2(new_n226), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n231), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(KEYINPUT80), .B(KEYINPUT39), .C1(new_n229), .C2(new_n231), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G57gat), .ZN(new_n246));
  INV_X1    g045(.A(G85gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n243), .A2(KEYINPUT39), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT40), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n239), .A3(new_n230), .A4(new_n241), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n231), .B1(new_n227), .B2(new_n228), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT77), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n255), .B2(KEYINPUT77), .ZN(new_n260));
  OR3_X1    g059(.A1(new_n259), .A2(new_n260), .A3(new_n250), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264));
  INV_X1    g063(.A(G64gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G183gat), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT24), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(KEYINPUT24), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT64), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR3_X1   g083(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n288), .B(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n279), .A2(new_n281), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT66), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n277), .A2(KEYINPUT25), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n295), .C1(new_n286), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT26), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT67), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n282), .C1(KEYINPUT26), .C2(new_n300), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT27), .B(G183gat), .Z(new_n304));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n304), .B2(G190gat), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n304), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n303), .A2(new_n274), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  AOI211_X1 g106(.A(KEYINPUT29), .B(new_n270), .C1(new_n297), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n297), .A2(new_n270), .A3(new_n307), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT73), .B(G218gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT22), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G211gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(KEYINPUT22), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n308), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n317), .B(G218gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n297), .A2(new_n307), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n269), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n268), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n308), .B2(new_n310), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n321), .A3(new_n309), .ZN(new_n328));
  INV_X1    g127(.A(new_n268), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(KEYINPUT30), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n327), .A2(new_n328), .A3(new_n332), .A4(new_n329), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n252), .A2(new_n253), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n263), .A2(new_n331), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G78gat), .B(G106gat), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT31), .ZN(new_n337));
  INV_X1    g136(.A(G50gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n323), .B1(new_n217), .B2(new_n236), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n321), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n319), .A2(new_n323), .A3(new_n217), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n217), .A2(new_n236), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G228gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n342), .A2(new_n343), .A3(new_n235), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n340), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT79), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n350), .A3(new_n340), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G22gat), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(new_n355), .A3(new_n350), .A4(new_n340), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n250), .B1(new_n259), .B2(new_n260), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n250), .C1(new_n259), .C2(new_n260), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n261), .A4(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n261), .A2(new_n362), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n328), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n327), .A2(KEYINPUT81), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n327), .A2(new_n328), .A3(new_n368), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n268), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n365), .B(new_n366), .C1(new_n370), .C2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT37), .B1(new_n320), .B2(new_n325), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n376), .A2(new_n268), .A3(new_n371), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n330), .B1(new_n377), .B2(new_n373), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n335), .B(new_n359), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT36), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n297), .A2(new_n226), .A3(new_n307), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n226), .B1(new_n297), .B2(new_n307), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n383), .A2(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT34), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n226), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n322), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n297), .A2(new_n226), .A3(new_n307), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(KEYINPUT72), .A3(new_n381), .A4(new_n382), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G71gat), .ZN(new_n400));
  INV_X1    g199(.A(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n389), .A3(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(KEYINPUT32), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT32), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n388), .B2(new_n389), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n402), .A2(KEYINPUT70), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT33), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n402), .A2(new_n405), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n398), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n403), .A2(KEYINPUT32), .A3(new_n410), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n388), .A2(new_n389), .B1(new_n406), .B2(KEYINPUT33), .ZN(new_n414));
  INV_X1    g213(.A(new_n402), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(new_n396), .A3(new_n397), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n380), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n390), .A3(new_n387), .A4(new_n395), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n396), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT36), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n365), .A2(new_n366), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n331), .A2(new_n333), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n359), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n379), .A2(new_n422), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n359), .A2(new_n412), .A3(new_n417), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT35), .B1(new_n429), .B2(new_n425), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n365), .A2(new_n366), .B1(new_n331), .B2(new_n333), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n419), .A2(new_n420), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT35), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n359), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G57gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(G64gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n265), .A2(G57gat), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT9), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G71gat), .A2(G78gat), .ZN(new_n441));
  OR2_X1    g240(.A1(G71gat), .A2(G78gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT9), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n265), .B2(G57gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n437), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(new_n438), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT21), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G15gat), .B(G22gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT16), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(G1gat), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(KEYINPUT88), .C1(G1gat), .C2(new_n457), .ZN(new_n460));
  INV_X1    g259(.A(G8gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n443), .A2(KEYINPUT21), .A3(new_n450), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G183gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n271), .A3(new_n463), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(G231gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n468), .ZN(new_n472));
  XNOR2_X1  g271(.A(G127gat), .B(G155gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(new_n315), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n470), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n470), .B2(new_n472), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n456), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n472), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n455), .A3(new_n476), .ZN(new_n482));
  AND2_X1   g281(.A1(G232gat), .A2(G233gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(KEYINPUT41), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT93), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(new_n272), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G218gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n338), .A2(G43gat), .ZN(new_n489));
  INV_X1    g288(.A(G43gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G50gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT15), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT14), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(new_n492), .ZN(new_n504));
  OR2_X1    g303(.A1(KEYINPUT86), .A2(G29gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT86), .A2(G29gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(G36gat), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n496), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT84), .B1(new_n489), .B2(new_n491), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n509), .A2(new_n510), .A3(new_n503), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n500), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT14), .B1(new_n497), .B2(new_n498), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n507), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n511), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n508), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  AOI22_X1  g323(.A1(KEYINPUT8), .A2(new_n524), .B1(new_n247), .B2(new_n267), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n247), .B2(new_n267), .ZN(new_n527));
  NAND3_X1  g326(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G99gat), .B(G106gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT17), .B(new_n508), .C1(new_n519), .C2(new_n520), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G134gat), .B(G162gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n531), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n521), .A2(new_n536), .B1(KEYINPUT41), .B2(new_n483), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n533), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n488), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n539), .A2(new_n488), .A3(new_n540), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n479), .A2(new_n482), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n545), .B(KEYINPUT10), .C1(new_n531), .C2(new_n451), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n451), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n529), .A2(new_n530), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n530), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n549), .A2(new_n443), .A3(new_n450), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT10), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT95), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n545), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n547), .A4(new_n546), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n547), .B2(new_n551), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(new_n299), .ZN(new_n565));
  INV_X1    g364(.A(G204gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570));
  INV_X1    g369(.A(new_n560), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n548), .A2(new_n571), .A3(new_n552), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n567), .B1(new_n572), .B2(new_n562), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n569), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G169gat), .B(G197gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT12), .Z(new_n583));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n496), .A2(new_n504), .A3(new_n507), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n516), .A2(new_n507), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT85), .B1(new_n499), .B2(new_n501), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT87), .B1(new_n588), .B2(new_n496), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n591), .B2(new_n462), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n460), .B(G8gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n521), .A2(KEYINPUT89), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n523), .A2(new_n462), .A3(new_n532), .ZN(new_n596));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n583), .B1(new_n600), .B2(KEYINPUT91), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n593), .B1(new_n591), .B2(KEYINPUT17), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n592), .A2(new_n594), .B1(new_n602), .B2(new_n523), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT18), .B1(new_n603), .B2(new_n597), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT18), .A4(new_n597), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n462), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n591), .A2(new_n462), .A3(new_n584), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT89), .B1(new_n521), .B2(new_n593), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n597), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n601), .A2(new_n606), .A3(new_n607), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n607), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT90), .B(new_n583), .C1(new_n616), .C2(new_n604), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n607), .A3(new_n614), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT90), .B1(new_n619), .B2(new_n583), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n577), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n436), .A2(new_n544), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n423), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G1gat), .ZN(G1324gat));
  INV_X1    g426(.A(new_n424), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n461), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n458), .A2(new_n461), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n624), .A2(new_n628), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT42), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT98), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(G1325gat));
  AOI21_X1  g439(.A(G15gat), .B1(new_n624), .B2(new_n432), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  INV_X1    g441(.A(new_n422), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(G15gat), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n624), .B2(new_n644), .ZN(G1326gat));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n426), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT43), .B(G22gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n543), .A2(new_n541), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n428), .B2(new_n435), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n479), .A2(new_n482), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n650), .A2(new_n651), .A3(new_n623), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n505), .A2(new_n506), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n625), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT45), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n652), .A2(new_n656), .A3(new_n625), .A4(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n622), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(new_n541), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n542), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n436), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n663), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n428), .B2(new_n435), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n662), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n674));
  INV_X1    g473(.A(new_n672), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n663), .B2(new_n650), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n662), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n423), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n658), .B1(new_n679), .B2(new_n653), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n658), .B(new_n682), .C1(new_n679), .C2(new_n653), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1328gat));
  NAND3_X1  g483(.A1(new_n652), .A2(new_n498), .A3(new_n628), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT46), .Z(new_n686));
  AOI21_X1  g485(.A(new_n424), .B1(new_n674), .B2(new_n678), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n498), .B2(new_n687), .ZN(G1329gat));
  OAI21_X1  g487(.A(G43gat), .B1(new_n673), .B2(new_n422), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n652), .A2(new_n490), .A3(new_n432), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(KEYINPUT47), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n678), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n643), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(G43gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n695), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g495(.A(G50gat), .B1(new_n673), .B2(new_n359), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n652), .A2(new_n338), .A3(new_n426), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(KEYINPUT48), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n698), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n693), .A2(new_n426), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(G50gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(G1331gat));
  NAND2_X1  g503(.A1(new_n619), .A2(new_n583), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n617), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n544), .A2(new_n615), .A3(new_n708), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n577), .B(new_n709), .C1(new_n428), .C2(new_n435), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n625), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT105), .B(G57gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n424), .B(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT49), .B(G64gat), .Z(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(G1333gat));
  NAND2_X1  g519(.A1(new_n710), .A2(new_n643), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G71gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n432), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(G71gat), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n426), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  INV_X1    g526(.A(new_n621), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n676), .A2(new_n651), .A3(new_n576), .A4(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729), .B2(new_n423), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n436), .A2(new_n651), .A3(new_n665), .A4(new_n728), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n247), .A4(new_n576), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n730), .B1(new_n736), .B2(new_n423), .ZN(G1336gat));
  OAI21_X1  g536(.A(G92gat), .B1(new_n729), .B2(new_n715), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n733), .A2(new_n267), .A3(new_n576), .A4(new_n716), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G92gat), .B1(new_n729), .B2(new_n424), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n739), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(new_n740), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n729), .B2(new_n422), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n734), .A2(new_n735), .A3(new_n401), .A4(new_n432), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n577), .ZN(G1338gat));
  OAI21_X1  g546(.A(G106gat), .B1(new_n729), .B2(new_n359), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n359), .A2(G106gat), .A3(new_n577), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT53), .B1(new_n733), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n733), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n748), .A2(new_n751), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n753), .A2(new_n758), .A3(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(new_n670), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n548), .A2(new_n552), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n561), .B(KEYINPUT54), .C1(new_n560), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n568), .B1(new_n572), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(KEYINPUT55), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n571), .B1(new_n553), .B2(new_n558), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n763), .A2(new_n560), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(new_n765), .ZN(new_n771));
  INV_X1    g570(.A(new_n766), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n773), .A3(new_n569), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n708), .B2(new_n615), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n616), .B1(new_n605), .B2(new_n604), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n603), .B2(new_n597), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n595), .A2(new_n596), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n779), .A2(KEYINPUT110), .A3(G229gat), .A4(G233gat), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT111), .B1(new_n611), .B2(new_n613), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n595), .A2(new_n782), .A3(new_n608), .A4(new_n612), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n778), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n776), .A2(new_n601), .B1(new_n784), .B2(new_n582), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n576), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n762), .B1(new_n775), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n582), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n615), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n774), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n670), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n661), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n709), .A2(new_n576), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n625), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(new_n359), .A3(new_n432), .A4(new_n715), .ZN(new_n797));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797), .B2(new_n728), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT112), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n429), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n715), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n728), .A2(G113gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n797), .B2(new_n577), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n801), .A2(G120gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n577), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807));
  INV_X1    g606(.A(new_n661), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n797), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n801), .ZN(new_n810));
  INV_X1    g609(.A(new_n651), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT113), .Z(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n628), .A2(new_n649), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT56), .Z(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n797), .B2(new_n649), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n426), .C1(new_n793), .C2(new_n794), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n771), .B2(new_n772), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n767), .A2(new_n569), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n621), .A2(new_n825), .B1(new_n785), .B2(new_n576), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n792), .B1(new_n826), .B2(new_n665), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n794), .B1(new_n827), .B2(new_n651), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT57), .B1(new_n828), .B2(new_n359), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n643), .A2(new_n716), .A3(new_n423), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G141gat), .B1(new_n831), .B2(new_n728), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n643), .A2(new_n359), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT116), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n795), .A2(KEYINPUT115), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n715), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n728), .A2(G141gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT58), .ZN(G1344gat));
  AND2_X1   g639(.A1(new_n835), .A2(new_n836), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n577), .A2(G148gat), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(new_n715), .A3(new_n834), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n621), .A2(new_n825), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n665), .B1(new_n846), .B2(new_n786), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n790), .A2(new_n774), .A3(new_n649), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n848), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(KEYINPUT120), .C1(new_n826), .C2(new_n665), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n651), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n794), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n359), .A2(KEYINPUT57), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n793), .A2(new_n794), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n359), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n860), .A2(new_n576), .A3(new_n830), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n844), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n822), .A2(new_n829), .A3(new_n830), .A4(new_n576), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n866), .A3(G148gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT117), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(new_n869), .A3(new_n866), .A4(G148gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n843), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT122), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n874), .B(new_n843), .C1(new_n864), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1345gat));
  OAI21_X1  g675(.A(new_n209), .B1(new_n837), .B2(new_n651), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n831), .A2(new_n209), .A3(new_n808), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT123), .ZN(G1346gat));
  NAND4_X1  g679(.A1(new_n841), .A2(new_n210), .A3(new_n816), .A4(new_n834), .ZN(new_n881));
  OAI21_X1  g680(.A(G162gat), .B1(new_n831), .B2(new_n762), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n861), .A2(new_n625), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n884), .A2(new_n628), .A3(new_n359), .A4(new_n432), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n728), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n861), .A2(new_n625), .A3(new_n715), .ZN(new_n887));
  INV_X1    g686(.A(new_n429), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(KEYINPUT124), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n621), .A2(new_n298), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(G1348gat));
  NOR3_X1   g694(.A1(new_n885), .A2(new_n299), .A3(new_n577), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n576), .A3(new_n892), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n299), .ZN(G1349gat));
  OAI21_X1  g697(.A(G183gat), .B1(new_n885), .B2(new_n808), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n651), .A2(new_n304), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n899), .B(KEYINPUT125), .C1(new_n889), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n885), .B2(new_n649), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(KEYINPUT61), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n670), .A2(new_n272), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n904), .A2(new_n905), .B1(new_n893), .B2(new_n906), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n643), .A2(new_n625), .A3(new_n424), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n860), .A2(new_n862), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n728), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n833), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n728), .A2(G197gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1352gat));
  INV_X1    g712(.A(new_n911), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n577), .B1(new_n915), .B2(KEYINPUT62), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n566), .A3(new_n916), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n917), .A2(new_n915), .A3(KEYINPUT62), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n915), .B2(KEYINPUT62), .ZN(new_n919));
  AND4_X1   g718(.A1(new_n576), .A2(new_n860), .A3(new_n862), .A4(new_n908), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n918), .B(new_n919), .C1(new_n566), .C2(new_n920), .ZN(G1353gat));
  OAI21_X1  g720(.A(G211gat), .B1(new_n909), .B2(new_n651), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT63), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n911), .A2(G211gat), .A3(new_n651), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT127), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(G1354gat));
  INV_X1    g726(.A(new_n312), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n909), .A2(new_n928), .A3(new_n649), .ZN(new_n929));
  AOI21_X1  g728(.A(G218gat), .B1(new_n914), .B2(new_n670), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1355gat));
endmodule


