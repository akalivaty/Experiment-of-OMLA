//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n452), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n468));
  INV_X1    g043(.A(G113), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G113), .A3(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(G2105), .B2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n460), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n478), .A2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n461), .B2(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n479), .A2(new_n480), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(new_n494), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n492), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n501), .A2(KEYINPUT69), .A3(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n516), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT70), .B(G51), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n513), .A2(new_n525), .ZN(new_n526));
  AND4_X1   g101(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n509), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n513), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n509), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n507), .A2(G81), .A3(new_n515), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n513), .A2(G43), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n535), .B(KEYINPUT72), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n554), .B2(new_n509), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n557));
  AND3_X1   g132(.A1(new_n501), .A2(KEYINPUT69), .A3(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(KEYINPUT69), .B1(new_n501), .B2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .A3(G651), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n555), .A2(new_n563), .B1(G91), .B2(new_n520), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n513), .A2(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n513), .B(G53), .C1(new_n566), .C2(new_n567), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n564), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  NAND4_X1  g152(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n526), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND3_X1  g154(.A1(new_n507), .A2(G87), .A3(new_n515), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n513), .A2(G49), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n560), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n583), .B1(new_n585), .B2(G651), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n583), .B(G651), .C1(new_n507), .C2(G74), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n582), .B1(new_n586), .B2(new_n588), .ZN(G288));
  OAI211_X1 g164(.A(G61), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n509), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n505), .A2(new_n506), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n593), .A2(G86), .A3(new_n557), .A4(new_n515), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n513), .A2(G48), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n592), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n560), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n509), .B1(new_n600), .B2(KEYINPUT78), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(KEYINPUT78), .B2(new_n600), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT79), .B(G85), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n520), .A2(new_n603), .B1(G47), .B2(new_n513), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(G290));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G301), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n507), .A2(G92), .A3(new_n515), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n507), .A2(KEYINPUT81), .A3(G92), .A4(new_n515), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n513), .A2(G54), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n509), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n613), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n610), .A2(new_n611), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n614), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n614), .A2(KEYINPUT82), .A3(new_n620), .A4(new_n618), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n607), .B1(new_n625), .B2(new_n606), .ZN(G284));
  AOI21_X1  g201(.A(new_n607), .B1(new_n625), .B2(new_n606), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G299), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n545), .A2(new_n606), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n632), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n634), .B1(new_n636), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n497), .A2(new_n465), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n483), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n481), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n460), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(KEYINPUT15), .B(G2435), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(G2072), .A2(G2078), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n442), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n675), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(KEYINPUT17), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n676), .C1(new_n673), .C2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n676), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2096), .B(G2100), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(new_n700), .B(new_n699), .S(new_n692), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(G229));
  XOR2_X1   g285(.A(KEYINPUT87), .B(G29), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n483), .A2(G131), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n481), .A2(G119), .ZN(new_n715));
  OR2_X1    g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT88), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(KEYINPUT88), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G24), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n730));
  XNOR2_X1  g305(.A(G290), .B(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n731), .B2(new_n726), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G1986), .ZN(new_n733));
  INV_X1    g308(.A(G1986), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(new_n729), .C1(new_n731), .C2(new_n726), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n722), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n592), .A2(new_n596), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G6), .B2(G16), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT32), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(KEYINPUT32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G1981), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n742), .A2(G1981), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n727), .A2(G22), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G166), .B2(new_n727), .ZN(new_n750));
  INV_X1    g325(.A(G1971), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n723), .A2(G23), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n580), .A2(new_n581), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n585), .A2(G651), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT77), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n754), .B1(new_n756), .B2(new_n587), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n753), .B1(new_n757), .B2(new_n723), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT33), .B(G1976), .Z(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n752), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n738), .B1(new_n748), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n764));
  INV_X1    g339(.A(new_n762), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n765), .A2(new_n737), .A3(new_n746), .A4(new_n747), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n736), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n736), .A2(new_n766), .A3(new_n763), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n768), .B(KEYINPUT36), .C1(KEYINPUT91), .C2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(KEYINPUT91), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  OR3_X1    g349(.A1(new_n712), .A2(KEYINPUT96), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT96), .B1(new_n712), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n773), .A2(G34), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G160), .ZN(new_n779));
  INV_X1    g354(.A(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2084), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT31), .B(G11), .Z(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G162), .A2(new_n712), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G35), .B2(new_n712), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT29), .B(G2090), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n787), .B1(new_n649), .B2(new_n711), .C1(new_n789), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n711), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n483), .A2(G140), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n481), .A2(G128), .ZN(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n780), .A2(G33), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G139), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n484), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n497), .A2(G127), .ZN(new_n810));
  INV_X1    g385(.A(G115), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n464), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(G2105), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n804), .B1(new_n815), .B2(G29), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(G2072), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(G2072), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n782), .B(new_n803), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n723), .A2(G21), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G168), .B2(new_n723), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT97), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n780), .A2(G32), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n465), .A2(G105), .ZN(new_n825));
  INV_X1    g400(.A(G141), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n484), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n481), .A2(G129), .ZN(new_n828));
  NAND3_X1  g403(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT26), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n824), .B1(new_n833), .B2(G29), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT27), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G1996), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n822), .A2(G1966), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n711), .A2(G27), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT99), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n496), .A2(new_n499), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n488), .A2(new_n491), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n843), .B1(new_n846), .B2(new_n712), .ZN(new_n847));
  INV_X1    g422(.A(G2078), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n789), .A2(new_n791), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n723), .A2(G5), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G171), .B2(new_n723), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(G1961), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n847), .A2(new_n848), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(G1961), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n849), .A2(new_n852), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n819), .A2(new_n841), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n822), .A2(G1966), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT98), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n727), .A2(G19), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n546), .B2(new_n727), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(G1341), .Z(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n726), .A2(G20), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT100), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT23), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G299), .B2(G16), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G1956), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT93), .ZN(new_n869));
  OR3_X1    g444(.A1(new_n869), .A2(G4), .A3(G16), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(G4), .B2(G16), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n623), .A2(new_n624), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n723), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT94), .B(G1348), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n862), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n770), .A2(new_n772), .A3(new_n876), .ZN(G311));
  NAND3_X1  g452(.A1(new_n770), .A2(new_n876), .A3(new_n772), .ZN(G150));
  NAND2_X1  g453(.A1(new_n625), .A2(G559), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n509), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n513), .A2(G55), .ZN(new_n884));
  INV_X1    g459(.A(G93), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n516), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n545), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n541), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n881), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  AOI21_X1  g469(.A(G860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(G860), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT37), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G145));
  XNOR2_X1  g474(.A(G164), .B(new_n799), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n815), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n833), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n815), .A2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n833), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n815), .A2(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n718), .B(KEYINPUT104), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n908), .A2(new_n640), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n640), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n483), .A2(G142), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n481), .A2(G130), .ZN(new_n912));
  OR2_X1    g487(.A1(G106), .A2(G2105), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n913), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n909), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n909), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(G160), .B(KEYINPUT103), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n649), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(G162), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n902), .A2(new_n918), .A3(new_n906), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G37), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n918), .B1(new_n902), .B2(new_n906), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(KEYINPUT105), .B2(new_n924), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n907), .A2(KEYINPUT105), .A3(new_n919), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n928), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n927), .A2(new_n933), .A3(KEYINPUT40), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT40), .B1(new_n927), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(G395));
  NAND2_X1  g511(.A1(new_n636), .A2(new_n892), .ZN(new_n937));
  NOR2_X1   g512(.A1(G299), .A2(new_n621), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G299), .A2(new_n621), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n887), .B1(new_n543), .B2(new_n544), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n890), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n635), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n937), .A2(new_n945), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n939), .B2(new_n940), .ZN(new_n949));
  INV_X1    g524(.A(new_n940), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n950), .A2(new_n938), .A3(KEYINPUT41), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT106), .B(new_n946), .C1(new_n947), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n757), .A2(new_n602), .A3(new_n604), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n757), .B1(new_n602), .B2(new_n604), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G290), .A2(G288), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT108), .A3(new_n955), .ZN(new_n960));
  XNOR2_X1  g535(.A(G166), .B(G305), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(new_n959), .A3(KEYINPUT108), .A4(new_n955), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT42), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n953), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n953), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g545(.A(G868), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n888), .A2(new_n606), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(G295));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n972), .ZN(G331));
  XNOR2_X1  g549(.A(G286), .B(G171), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n892), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n943), .A2(new_n975), .A3(new_n890), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n978), .C1(new_n949), .C2(new_n951), .ZN(new_n979));
  INV_X1    g554(.A(new_n965), .ZN(new_n980));
  INV_X1    g555(.A(new_n975), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n944), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n942), .B1(new_n982), .B2(new_n977), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n979), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n926), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n980), .B1(new_n979), .B2(new_n983), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT41), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n941), .A2(new_n988), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n950), .A2(new_n938), .A3(new_n948), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n976), .A4(new_n978), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n983), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n965), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n994), .A3(new_n926), .A4(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n926), .A3(new_n984), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(new_n986), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(new_n994), .A3(new_n926), .A4(new_n984), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1002), .A3(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(G397));
  AOI21_X1  g579(.A(G1384), .B1(new_n844), .B2(new_n845), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n470), .A2(new_n472), .ZN(new_n1011));
  INV_X1    g586(.A(G125), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n479), .B2(new_n480), .ZN(new_n1013));
  OAI21_X1  g588(.A(G2105), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n463), .A2(new_n466), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(G40), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1996), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT111), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1017), .B2(G1996), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n833), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n799), .B(G2067), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n833), .A2(G1996), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1017), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n718), .B(new_n721), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n602), .A2(new_n734), .A3(new_n604), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G290), .A2(G1986), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G166), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1016), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT112), .B(new_n1009), .C1(G164), .C2(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1014), .A2(new_n1015), .A3(G40), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n846), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2090), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n751), .A2(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1036), .B1(new_n1049), .B2(new_n1033), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n751), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n846), .A2(G160), .A3(G40), .A4(new_n1045), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  NAND4_X1  g633(.A1(G288), .A2(new_n1057), .A3(G8), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1033), .B1(new_n1043), .B2(new_n1005), .ZN(new_n1062));
  OAI211_X1 g637(.A(G1976), .B(new_n582), .C1(new_n586), .C2(new_n588), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT113), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT113), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G305), .A2(G1981), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT114), .B(G1981), .Z(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n739), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n592), .A2(new_n596), .A3(new_n1073), .A4(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1069), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT49), .B(new_n1069), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1062), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT117), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1068), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1056), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n1045), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(new_n1043), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(G2078), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT124), .B(G1961), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1087), .A2(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1041), .B2(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1086), .A2(new_n1043), .A3(new_n1089), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1096), .A2(new_n1097), .B1(new_n1010), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1090), .A2(KEYINPUT125), .A3(new_n1091), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(G301), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1085), .A2(new_n1043), .A3(new_n1086), .ZN(new_n1104));
  INV_X1    g679(.A(G1966), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1042), .A2(new_n1046), .A3(new_n1107), .A4(new_n1043), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(G168), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(G168), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(G8), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1102), .A2(new_n1103), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1098), .A2(new_n1010), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1093), .A2(new_n1116), .A3(new_n1100), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G171), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1092), .A2(new_n1093), .A3(G301), .ZN(new_n1120));
  AND4_X1   g695(.A1(KEYINPUT126), .A2(new_n1119), .A3(KEYINPUT54), .A4(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(KEYINPUT54), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT126), .B1(new_n1122), .B2(new_n1119), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1084), .B(new_n1115), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT56), .B(G2072), .Z(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT118), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1090), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT120), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(KEYINPUT119), .A3(new_n1040), .A4(new_n1126), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT57), .B1(new_n569), .B2(new_n570), .ZN(new_n1139));
  AOI22_X1  g714(.A1(G299), .A2(KEYINPUT57), .B1(new_n564), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1134), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n623), .B2(new_n624), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1057), .A2(G2067), .ZN(new_n1150));
  INV_X1    g725(.A(G1348), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1090), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n623), .A2(new_n1148), .A3(new_n624), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n625), .A2(KEYINPUT60), .A3(new_n1152), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1038), .A2(new_n1039), .A3(new_n837), .A4(new_n1040), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1057), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1057), .A2(KEYINPUT121), .A3(new_n1157), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1156), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1162), .A2(new_n546), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1162), .B2(new_n546), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1154), .A2(new_n1155), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1141), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1136), .A2(new_n1140), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT61), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1142), .A2(new_n1145), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1147), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1142), .B1(new_n872), .B2(new_n1152), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1169), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1124), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1095), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1112), .A2(new_n1114), .A3(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1084), .A2(new_n1179), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1080), .A2(new_n1055), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G288), .A2(G1976), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  OAI22_X1  g762(.A1(new_n1185), .A2(new_n1187), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1184), .B1(new_n1062), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1033), .B(G286), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n1084), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(KEYINPUT63), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1056), .A2(new_n1080), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1183), .B(new_n1189), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1032), .B1(new_n1177), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1017), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n719), .A2(new_n721), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1022), .A2(new_n1025), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n799), .A2(G2067), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1196), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT48), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1019), .A2(KEYINPUT46), .A3(new_n1021), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1017), .B1(new_n904), .B2(new_n1023), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1203), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g786(.A(KEYINPUT47), .B(new_n1209), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1212));
  OAI221_X1 g787(.A(new_n1200), .B1(new_n1028), .B2(new_n1202), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1195), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g790(.A1(new_n687), .A2(G319), .A3(new_n688), .ZN(new_n1217));
  XNOR2_X1  g791(.A(new_n1217), .B(KEYINPUT127), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n669), .B(new_n1218), .C1(new_n708), .C2(new_n709), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n933), .B2(new_n927), .ZN(new_n1220));
  AND2_X1   g794(.A1(new_n1220), .A2(new_n996), .ZN(G308));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n996), .ZN(G225));
endmodule


