

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724;

  XNOR2_X1 U367 ( .A(n468), .B(KEYINPUT105), .ZN(n555) );
  NOR2_X1 U368 ( .A1(n722), .A2(n724), .ZN(n495) );
  XNOR2_X1 U369 ( .A(n570), .B(n344), .ZN(n467) );
  AND2_X1 U370 ( .A1(n552), .A2(n438), .ZN(n570) );
  BUF_X1 U371 ( .A(n535), .Z(n345) );
  AND2_X1 U372 ( .A1(n537), .A2(n348), .ZN(n494) );
  INV_X1 U373 ( .A(n439), .ZN(n344) );
  XNOR2_X1 U374 ( .A(n416), .B(n415), .ZN(n510) );
  AND2_X1 U375 ( .A1(n482), .A2(n639), .ZN(n558) );
  OR2_X1 U376 ( .A1(n604), .A2(n405), .ZN(n411) );
  XNOR2_X1 U377 ( .A(n460), .B(n459), .ZN(n703) );
  XNOR2_X1 U378 ( .A(n351), .B(n346), .ZN(n460) );
  XNOR2_X1 U379 ( .A(n390), .B(n389), .ZN(n446) );
  XNOR2_X1 U380 ( .A(n455), .B(n347), .ZN(n346) );
  INV_X1 U381 ( .A(KEYINPUT23), .ZN(n347) );
  XNOR2_X1 U382 ( .A(G119), .B(G116), .ZN(n388) );
  INV_X1 U383 ( .A(G953), .ZN(n714) );
  NAND2_X1 U384 ( .A1(n586), .A2(n585), .ZN(n635) );
  NOR2_X2 U385 ( .A1(n515), .A2(n656), .ZN(n492) );
  XNOR2_X2 U386 ( .A(n490), .B(n489), .ZN(n515) );
  XNOR2_X2 U387 ( .A(n530), .B(n529), .ZN(n708) );
  NOR2_X1 U388 ( .A1(G953), .A2(G237), .ZN(n443) );
  INV_X1 U389 ( .A(G110), .ZN(n469) );
  OR2_X1 U390 ( .A1(n501), .A2(n655), .ZN(n531) );
  XNOR2_X1 U391 ( .A(G475), .B(n372), .ZN(n514) );
  AND2_X1 U392 ( .A1(n642), .A2(n548), .ZN(n639) );
  XNOR2_X1 U393 ( .A(n482), .B(KEYINPUT1), .ZN(n638) );
  NOR2_X4 U394 ( .A1(n635), .A2(n587), .ZN(n624) );
  BUF_X1 U395 ( .A(n692), .Z(n348) );
  XNOR2_X2 U396 ( .A(n540), .B(n539), .ZN(n665) );
  NOR2_X2 U397 ( .A1(n549), .A2(n561), .ZN(n540) );
  XNOR2_X1 U398 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U399 ( .A(KEYINPUT39), .ZN(n491) );
  INV_X1 U400 ( .A(KEYINPUT104), .ZN(n439) );
  XNOR2_X1 U401 ( .A(n429), .B(G137), .ZN(n430) );
  XNOR2_X1 U402 ( .A(n425), .B(n424), .ZN(n541) );
  XNOR2_X1 U403 ( .A(n528), .B(KEYINPUT79), .ZN(n529) );
  INV_X1 U404 ( .A(n458), .ZN(n368) );
  XNOR2_X1 U405 ( .A(n365), .B(n364), .ZN(n369) );
  XNOR2_X1 U406 ( .A(n359), .B(n358), .ZN(n365) );
  INV_X1 U407 ( .A(KEYINPUT33), .ZN(n539) );
  XOR2_X1 U408 ( .A(KEYINPUT97), .B(n514), .Z(n505) );
  BUF_X1 U409 ( .A(n541), .Z(n563) );
  NOR2_X1 U410 ( .A1(n532), .A2(n638), .ZN(n534) );
  NOR2_X1 U411 ( .A1(n512), .A2(n519), .ZN(n349) );
  AND2_X1 U412 ( .A1(n658), .A2(n642), .ZN(n350) );
  AND2_X1 U413 ( .A1(n456), .A2(G221), .ZN(n351) );
  AND2_X1 U414 ( .A1(n496), .A2(n466), .ZN(n352) );
  AND2_X1 U415 ( .A1(n477), .A2(n482), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n497), .B(KEYINPUT6), .ZN(n549) );
  OR2_X1 U417 ( .A1(n721), .A2(n554), .ZN(n556) );
  INV_X1 U418 ( .A(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U419 ( .A(G131), .B(KEYINPUT4), .ZN(n429) );
  INV_X1 U420 ( .A(n484), .ZN(n485) );
  XNOR2_X1 U421 ( .A(G140), .B(KEYINPUT10), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n366), .B(G125), .ZN(n399) );
  INV_X1 U423 ( .A(KEYINPUT19), .ZN(n415) );
  XNOR2_X1 U424 ( .A(n399), .B(n367), .ZN(n458) );
  INV_X1 U425 ( .A(KEYINPUT73), .ZN(n489) );
  AND2_X1 U426 ( .A1(n595), .A2(n701), .ZN(n709) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n588) );
  INV_X1 U428 ( .A(KEYINPUT43), .ZN(n533) );
  XNOR2_X1 U429 ( .A(n428), .B(n427), .ZN(n552) );
  XNOR2_X1 U430 ( .A(n493), .B(KEYINPUT101), .ZN(n692) );
  AND2_X1 U431 ( .A1(n591), .A2(G953), .ZN(n707) );
  XOR2_X1 U432 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n355) );
  XNOR2_X1 U433 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n354) );
  XNOR2_X1 U434 ( .A(n355), .B(n354), .ZN(n359) );
  XNOR2_X1 U435 ( .A(G131), .B(G143), .ZN(n357) );
  NAND2_X1 U436 ( .A1(G214), .A2(n443), .ZN(n361) );
  XNOR2_X1 U437 ( .A(G113), .B(G104), .ZN(n360) );
  XNOR2_X1 U438 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U439 ( .A(KEYINPUT95), .B(G122), .Z(n362) );
  XNOR2_X1 U440 ( .A(n363), .B(n362), .ZN(n364) );
  INV_X1 U441 ( .A(G146), .ZN(n366) );
  NOR2_X1 U442 ( .A1(G902), .A2(n588), .ZN(n371) );
  XNOR2_X1 U443 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U445 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n382) );
  XNOR2_X2 U446 ( .A(G143), .B(G128), .ZN(n400) );
  XNOR2_X1 U447 ( .A(n400), .B(G134), .ZN(n431) );
  XOR2_X1 U448 ( .A(KEYINPUT9), .B(G122), .Z(n374) );
  XNOR2_X1 U449 ( .A(G116), .B(G107), .ZN(n373) );
  XNOR2_X1 U450 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U451 ( .A(n431), .B(n375), .ZN(n380) );
  NAND2_X1 U452 ( .A1(G234), .A2(n714), .ZN(n376) );
  XOR2_X1 U453 ( .A(KEYINPUT8), .B(n376), .Z(n456) );
  NAND2_X1 U454 ( .A1(G217), .A2(n456), .ZN(n378) );
  XOR2_X1 U455 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n377) );
  XNOR2_X1 U456 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U457 ( .A(n380), .B(n379), .ZN(n626) );
  NOR2_X1 U458 ( .A1(G902), .A2(n626), .ZN(n381) );
  XNOR2_X1 U459 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U460 ( .A(G478), .B(n383), .ZN(n513) );
  NOR2_X1 U461 ( .A1(n514), .A2(n513), .ZN(n658) );
  XNOR2_X1 U462 ( .A(KEYINPUT15), .B(G902), .ZN(n587) );
  NAND2_X1 U463 ( .A1(n587), .A2(G234), .ZN(n385) );
  XNOR2_X1 U464 ( .A(KEYINPUT20), .B(KEYINPUT86), .ZN(n384) );
  XNOR2_X1 U465 ( .A(n385), .B(n384), .ZN(n461) );
  NAND2_X1 U466 ( .A1(n461), .A2(G221), .ZN(n386) );
  XOR2_X1 U467 ( .A(KEYINPUT88), .B(n386), .Z(n387) );
  XNOR2_X1 U468 ( .A(n387), .B(KEYINPUT21), .ZN(n642) );
  XNOR2_X1 U469 ( .A(n388), .B(KEYINPUT3), .ZN(n390) );
  XNOR2_X1 U470 ( .A(G113), .B(KEYINPUT66), .ZN(n389) );
  XNOR2_X1 U471 ( .A(KEYINPUT16), .B(G122), .ZN(n391) );
  XNOR2_X1 U472 ( .A(n446), .B(n391), .ZN(n395) );
  XNOR2_X1 U473 ( .A(G107), .B(G104), .ZN(n392) );
  XNOR2_X1 U474 ( .A(n392), .B(n469), .ZN(n394) );
  XNOR2_X1 U475 ( .A(G101), .B(KEYINPUT72), .ZN(n393) );
  XNOR2_X1 U476 ( .A(n394), .B(n393), .ZN(n435) );
  XNOR2_X1 U477 ( .A(n395), .B(n435), .ZN(n620) );
  XNOR2_X1 U478 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n397) );
  NAND2_X1 U479 ( .A1(n714), .A2(G224), .ZN(n396) );
  XNOR2_X1 U480 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U481 ( .A(n399), .B(n398), .ZN(n403) );
  XNOR2_X1 U482 ( .A(KEYINPUT80), .B(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U483 ( .A(n400), .B(n401), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U485 ( .A(n620), .B(n404), .ZN(n604) );
  INV_X1 U486 ( .A(n587), .ZN(n405) );
  INV_X1 U487 ( .A(G902), .ZN(n450) );
  INV_X1 U488 ( .A(G237), .ZN(n406) );
  NAND2_X1 U489 ( .A1(n450), .A2(n406), .ZN(n412) );
  NAND2_X1 U490 ( .A1(n412), .A2(G210), .ZN(n407) );
  XNOR2_X1 U491 ( .A(n407), .B(KEYINPUT83), .ZN(n409) );
  XNOR2_X1 U492 ( .A(KEYINPUT75), .B(KEYINPUT82), .ZN(n408) );
  XNOR2_X1 U493 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X2 U494 ( .A(n411), .B(n410), .ZN(n535) );
  NAND2_X1 U495 ( .A1(n412), .A2(G214), .ZN(n414) );
  INV_X1 U496 ( .A(KEYINPUT84), .ZN(n413) );
  XNOR2_X1 U497 ( .A(n414), .B(n413), .ZN(n655) );
  NOR2_X2 U498 ( .A1(n535), .A2(n655), .ZN(n416) );
  XOR2_X1 U499 ( .A(KEYINPUT14), .B(KEYINPUT85), .Z(n418) );
  NAND2_X1 U500 ( .A1(G234), .A2(G237), .ZN(n417) );
  XNOR2_X1 U501 ( .A(n418), .B(n417), .ZN(n419) );
  AND2_X1 U502 ( .A1(n419), .A2(G952), .ZN(n669) );
  AND2_X1 U503 ( .A1(n669), .A2(n714), .ZN(n473) );
  INV_X1 U504 ( .A(n473), .ZN(n421) );
  INV_X1 U505 ( .A(G898), .ZN(n616) );
  NAND2_X1 U506 ( .A1(G953), .A2(n616), .ZN(n621) );
  NAND2_X1 U507 ( .A1(G902), .A2(n419), .ZN(n470) );
  OR2_X1 U508 ( .A1(n621), .A2(n470), .ZN(n420) );
  NAND2_X1 U509 ( .A1(n421), .A2(n420), .ZN(n422) );
  NAND2_X1 U510 ( .A1(n510), .A2(n422), .ZN(n425) );
  INV_X1 U511 ( .A(KEYINPUT64), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n423), .B(KEYINPUT0), .ZN(n424) );
  NAND2_X1 U513 ( .A1(n350), .A2(n541), .ZN(n428) );
  XNOR2_X1 U514 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U515 ( .A(n426), .B(KEYINPUT68), .ZN(n427) );
  XNOR2_X1 U516 ( .A(n431), .B(n430), .ZN(n711) );
  XNOR2_X1 U517 ( .A(G146), .B(n711), .ZN(n449) );
  XOR2_X1 U518 ( .A(KEYINPUT74), .B(G140), .Z(n433) );
  NAND2_X1 U519 ( .A1(G227), .A2(n714), .ZN(n432) );
  XNOR2_X1 U520 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U521 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U522 ( .A(n449), .B(n436), .ZN(n631) );
  NAND2_X1 U523 ( .A1(n631), .A2(n450), .ZN(n437) );
  XNOR2_X1 U524 ( .A(n437), .B(G469), .ZN(n482) );
  INV_X1 U525 ( .A(n638), .ZN(n438) );
  XOR2_X1 U526 ( .A(G101), .B(KEYINPUT71), .Z(n442) );
  XNOR2_X1 U527 ( .A(KEYINPUT5), .B(KEYINPUT89), .ZN(n441) );
  XNOR2_X1 U528 ( .A(n442), .B(n441), .ZN(n445) );
  NAND2_X1 U529 ( .A1(n443), .A2(G210), .ZN(n444) );
  XNOR2_X1 U530 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U531 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U532 ( .A(n449), .B(n448), .ZN(n598) );
  NAND2_X1 U533 ( .A1(n598), .A2(n450), .ZN(n452) );
  XNOR2_X1 U534 ( .A(G472), .B(KEYINPUT67), .ZN(n451) );
  XNOR2_X2 U535 ( .A(n452), .B(n451), .ZN(n496) );
  XOR2_X1 U536 ( .A(G110), .B(G119), .Z(n454) );
  XNOR2_X1 U537 ( .A(G128), .B(G137), .ZN(n453) );
  XNOR2_X1 U538 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U539 ( .A(n458), .B(KEYINPUT24), .ZN(n459) );
  NOR2_X2 U540 ( .A1(G902), .A2(n703), .ZN(n465) );
  AND2_X1 U541 ( .A1(n461), .A2(G217), .ZN(n463) );
  XNOR2_X1 U542 ( .A(KEYINPUT25), .B(KEYINPUT87), .ZN(n462) );
  XNOR2_X1 U543 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X2 U544 ( .A(n465), .B(n464), .ZN(n548) );
  INV_X1 U545 ( .A(n548), .ZN(n466) );
  NAND2_X1 U546 ( .A1(n467), .A2(n352), .ZN(n468) );
  XNOR2_X1 U547 ( .A(n555), .B(n469), .ZN(G12) );
  XOR2_X1 U548 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n481) );
  OR2_X1 U549 ( .A1(n714), .A2(n470), .ZN(n471) );
  NOR2_X1 U550 ( .A1(G900), .A2(n471), .ZN(n472) );
  NOR2_X1 U551 ( .A1(n473), .A2(n472), .ZN(n484) );
  NOR2_X1 U552 ( .A1(n484), .A2(n548), .ZN(n474) );
  NAND2_X1 U553 ( .A1(n642), .A2(n474), .ZN(n498) );
  OR2_X1 U554 ( .A1(n498), .A2(n496), .ZN(n475) );
  XNOR2_X1 U555 ( .A(n475), .B(KEYINPUT28), .ZN(n476) );
  XNOR2_X1 U556 ( .A(KEYINPUT109), .B(n476), .ZN(n477) );
  INV_X1 U557 ( .A(KEYINPUT38), .ZN(n478) );
  XNOR2_X1 U558 ( .A(n535), .B(n478), .ZN(n656) );
  NOR2_X1 U559 ( .A1(n656), .A2(n655), .ZN(n661) );
  NAND2_X1 U560 ( .A1(n658), .A2(n661), .ZN(n479) );
  XNOR2_X1 U561 ( .A(KEYINPUT41), .B(n479), .ZN(n653) );
  NAND2_X1 U562 ( .A1(n353), .A2(n653), .ZN(n480) );
  XNOR2_X1 U563 ( .A(n481), .B(n480), .ZN(n722) );
  XNOR2_X1 U564 ( .A(KEYINPUT108), .B(n558), .ZN(n488) );
  NOR2_X1 U565 ( .A1(n496), .A2(n655), .ZN(n483) );
  XNOR2_X1 U566 ( .A(n483), .B(KEYINPUT30), .ZN(n486) );
  AND2_X1 U567 ( .A1(n486), .A2(n485), .ZN(n487) );
  NAND2_X1 U568 ( .A1(n488), .A2(n487), .ZN(n490) );
  XNOR2_X1 U569 ( .A(n492), .B(n491), .ZN(n537) );
  INV_X1 U570 ( .A(n513), .ZN(n506) );
  NAND2_X1 U571 ( .A1(n505), .A2(n506), .ZN(n493) );
  XNOR2_X1 U572 ( .A(n494), .B(KEYINPUT40), .ZN(n724) );
  XNOR2_X1 U573 ( .A(n495), .B(KEYINPUT46), .ZN(n504) );
  XOR2_X1 U574 ( .A(n496), .B(KEYINPUT102), .Z(n497) );
  NOR2_X1 U575 ( .A1(n549), .A2(n498), .ZN(n499) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(n499), .ZN(n500) );
  NAND2_X1 U577 ( .A1(n500), .A2(n348), .ZN(n501) );
  NOR2_X1 U578 ( .A1(n531), .A2(n345), .ZN(n502) );
  XNOR2_X1 U579 ( .A(n502), .B(KEYINPUT36), .ZN(n503) );
  NAND2_X1 U580 ( .A1(n503), .A2(n638), .ZN(n698) );
  AND2_X1 U581 ( .A1(n504), .A2(n698), .ZN(n527) );
  NOR2_X1 U582 ( .A1(n506), .A2(n505), .ZN(n694) );
  NOR2_X1 U583 ( .A1(n348), .A2(n694), .ZN(n659) );
  INV_X1 U584 ( .A(KEYINPUT47), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(KEYINPUT65), .ZN(n507) );
  NOR2_X1 U586 ( .A1(n659), .A2(n507), .ZN(n508) );
  XNOR2_X1 U587 ( .A(n508), .B(KEYINPUT70), .ZN(n509) );
  NOR2_X1 U588 ( .A1(KEYINPUT77), .A2(n509), .ZN(n512) );
  BUF_X1 U589 ( .A(n510), .Z(n511) );
  NAND2_X1 U590 ( .A1(n353), .A2(n511), .ZN(n519) );
  AND2_X1 U591 ( .A1(n514), .A2(n513), .ZN(n544) );
  INV_X1 U592 ( .A(n515), .ZN(n516) );
  NAND2_X1 U593 ( .A1(n544), .A2(n516), .ZN(n517) );
  OR2_X1 U594 ( .A1(n345), .A2(n517), .ZN(n689) );
  NAND2_X1 U595 ( .A1(KEYINPUT77), .A2(n522), .ZN(n518) );
  NAND2_X1 U596 ( .A1(n689), .A2(n518), .ZN(n524) );
  INV_X1 U597 ( .A(n519), .ZN(n690) );
  NOR2_X1 U598 ( .A1(n690), .A2(KEYINPUT77), .ZN(n520) );
  NOR2_X1 U599 ( .A1(n659), .A2(n520), .ZN(n521) );
  NOR2_X1 U600 ( .A1(n522), .A2(n521), .ZN(n523) );
  OR2_X1 U601 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U602 ( .A1(n349), .A2(n525), .ZN(n526) );
  NAND2_X1 U603 ( .A1(n527), .A2(n526), .ZN(n530) );
  INV_X1 U604 ( .A(KEYINPUT48), .ZN(n528) );
  XOR2_X1 U605 ( .A(KEYINPUT107), .B(n531), .Z(n532) );
  XNOR2_X1 U606 ( .A(n534), .B(n533), .ZN(n536) );
  NAND2_X1 U607 ( .A1(n536), .A2(n345), .ZN(n595) );
  NAND2_X1 U608 ( .A1(n537), .A2(n694), .ZN(n701) );
  NAND2_X1 U609 ( .A1(n709), .A2(KEYINPUT76), .ZN(n538) );
  NOR2_X1 U610 ( .A1(n708), .A2(n538), .ZN(n575) );
  NAND2_X1 U611 ( .A1(n639), .A2(n638), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n665), .A2(n563), .ZN(n543) );
  INV_X1 U613 ( .A(KEYINPUT34), .ZN(n542) );
  XNOR2_X1 U614 ( .A(n543), .B(n542), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n546), .B(KEYINPUT35), .ZN(n721) );
  INV_X1 U617 ( .A(KEYINPUT103), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n548), .B(n547), .ZN(n641) );
  INV_X1 U619 ( .A(n549), .ZN(n568) );
  NOR2_X1 U620 ( .A1(n641), .A2(n568), .ZN(n550) );
  AND2_X1 U621 ( .A1(n638), .A2(n550), .ZN(n551) );
  NAND2_X1 U622 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n553), .B(KEYINPUT32), .ZN(n723) );
  INV_X1 U624 ( .A(n723), .ZN(n554) );
  NOR2_X2 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n557), .B(KEYINPUT44), .ZN(n573) );
  AND2_X1 U627 ( .A1(n558), .A2(n496), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n559), .A2(n563), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT90), .B(n560), .Z(n682) );
  OR2_X1 U630 ( .A1(n496), .A2(n561), .ZN(n650) );
  INV_X1 U631 ( .A(n650), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT31), .B(KEYINPUT91), .Z(n564) );
  XNOR2_X1 U634 ( .A(n565), .B(n564), .ZN(n695) );
  NOR2_X1 U635 ( .A1(n682), .A2(n695), .ZN(n566) );
  NOR2_X1 U636 ( .A1(n566), .A2(n659), .ZN(n571) );
  INV_X1 U637 ( .A(n641), .ZN(n567) );
  NOR2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n677) );
  NOR2_X1 U640 ( .A1(n571), .A2(n677), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X2 U642 ( .A(n574), .B(KEYINPUT45), .ZN(n611) );
  NAND2_X1 U643 ( .A1(n575), .A2(n611), .ZN(n577) );
  INV_X1 U644 ( .A(KEYINPUT2), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n701), .A2(KEYINPUT2), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n578), .A2(KEYINPUT76), .ZN(n581) );
  INV_X1 U648 ( .A(KEYINPUT76), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n579), .A2(n701), .ZN(n580) );
  AND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n595), .A2(n582), .ZN(n583) );
  NOR2_X1 U652 ( .A1(n708), .A2(n583), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n584), .A2(n611), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n624), .A2(G475), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT59), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n592) );
  INV_X1 U657 ( .A(G952), .ZN(n591) );
  INV_X1 U658 ( .A(n707), .ZN(n607) );
  NAND2_X1 U659 ( .A1(n592), .A2(n607), .ZN(n594) );
  INV_X1 U660 ( .A(KEYINPUT60), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n594), .B(n593), .ZN(G60) );
  XNOR2_X1 U662 ( .A(n595), .B(G140), .ZN(G42) );
  NAND2_X1 U663 ( .A1(n624), .A2(G472), .ZN(n600) );
  XNOR2_X1 U664 ( .A(KEYINPUT81), .B(KEYINPUT111), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT62), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n600), .B(n599), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n601), .A2(n607), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U670 ( .A1(n624), .A2(G210), .ZN(n606) );
  XNOR2_X1 U671 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n608), .A2(n607), .ZN(n610) );
  XOR2_X1 U675 ( .A(KEYINPUT78), .B(KEYINPUT56), .Z(n609) );
  XNOR2_X1 U676 ( .A(n610), .B(n609), .ZN(G51) );
  BUF_X1 U677 ( .A(n611), .Z(n612) );
  NAND2_X1 U678 ( .A1(n612), .A2(n714), .ZN(n613) );
  XOR2_X1 U679 ( .A(n613), .B(KEYINPUT126), .Z(n619) );
  NAND2_X1 U680 ( .A1(G953), .A2(G224), .ZN(n614) );
  XOR2_X1 U681 ( .A(KEYINPUT61), .B(n614), .Z(n615) );
  NOR2_X1 U682 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U683 ( .A(KEYINPUT125), .B(n617), .Z(n618) );
  NOR2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U685 ( .A1(n620), .A2(n621), .ZN(n622) );
  XNOR2_X1 U686 ( .A(n623), .B(n622), .ZN(G69) );
  BUF_X2 U687 ( .A(n624), .Z(n702) );
  NAND2_X1 U688 ( .A1(n702), .A2(G478), .ZN(n628) );
  XOR2_X1 U689 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n625) );
  XNOR2_X1 U690 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U691 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U692 ( .A1(n629), .A2(n707), .ZN(G63) );
  NAND2_X1 U693 ( .A1(n702), .A2(G469), .ZN(n633) );
  XNOR2_X1 U694 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n630) );
  XNOR2_X1 U695 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U696 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X1 U697 ( .A1(n634), .A2(n707), .ZN(G54) );
  BUF_X1 U698 ( .A(n635), .Z(n674) );
  NAND2_X1 U699 ( .A1(n665), .A2(n653), .ZN(n636) );
  XOR2_X1 U700 ( .A(KEYINPUT120), .B(n636), .Z(n637) );
  NOR2_X1 U701 ( .A1(n637), .A2(G953), .ZN(n672) );
  NOR2_X1 U702 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U703 ( .A(KEYINPUT50), .B(n640), .Z(n648) );
  INV_X1 U704 ( .A(n496), .ZN(n645) );
  NOR2_X1 U705 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U706 ( .A(KEYINPUT49), .B(n643), .Z(n644) );
  NOR2_X1 U707 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U708 ( .A(KEYINPUT118), .B(n646), .ZN(n647) );
  NAND2_X1 U709 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U710 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U711 ( .A(KEYINPUT51), .B(n651), .Z(n652) );
  NAND2_X1 U712 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U713 ( .A(KEYINPUT119), .B(n654), .Z(n667) );
  NAND2_X1 U714 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U715 ( .A1(n658), .A2(n657), .ZN(n663) );
  INV_X1 U716 ( .A(n659), .ZN(n660) );
  NAND2_X1 U717 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U718 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U719 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U720 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U721 ( .A(n668), .B(KEYINPUT52), .ZN(n670) );
  NAND2_X1 U722 ( .A1(n670), .A2(n669), .ZN(n671) );
  AND2_X1 U723 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U724 ( .A1(n674), .A2(n673), .ZN(n676) );
  XNOR2_X1 U725 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n675) );
  XNOR2_X1 U726 ( .A(n676), .B(n675), .ZN(G75) );
  XOR2_X1 U727 ( .A(G101), .B(n677), .Z(G3) );
  NAND2_X1 U728 ( .A1(n682), .A2(n348), .ZN(n678) );
  XNOR2_X1 U729 ( .A(n678), .B(KEYINPUT112), .ZN(n679) );
  XNOR2_X1 U730 ( .A(G104), .B(n679), .ZN(G6) );
  XOR2_X1 U731 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n681) );
  XNOR2_X1 U732 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U733 ( .A(n681), .B(n680), .ZN(n686) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT26), .ZN(n684) );
  NAND2_X1 U735 ( .A1(n694), .A2(n682), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U737 ( .A(n686), .B(n685), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U739 ( .A1(n690), .A2(n694), .ZN(n687) );
  XNOR2_X1 U740 ( .A(n688), .B(n687), .ZN(G30) );
  XNOR2_X1 U741 ( .A(G143), .B(n689), .ZN(G45) );
  NAND2_X1 U742 ( .A1(n690), .A2(n348), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n691), .B(G146), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n695), .A2(n348), .ZN(n693) );
  XNOR2_X1 U745 ( .A(n693), .B(G113), .ZN(G15) );
  NAND2_X1 U746 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U747 ( .A(n696), .B(KEYINPUT116), .ZN(n697) );
  XNOR2_X1 U748 ( .A(G116), .B(n697), .ZN(G18) );
  XNOR2_X1 U749 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U751 ( .A(G125), .B(n700), .ZN(G27) );
  XNOR2_X1 U752 ( .A(G134), .B(n701), .ZN(G36) );
  NAND2_X1 U753 ( .A1(n702), .A2(G217), .ZN(n705) );
  XNOR2_X1 U754 ( .A(n703), .B(KEYINPUT124), .ZN(n704) );
  XNOR2_X1 U755 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U756 ( .A1(n707), .A2(n706), .ZN(G66) );
  INV_X1 U757 ( .A(n708), .ZN(n710) );
  NAND2_X1 U758 ( .A1(n710), .A2(n709), .ZN(n713) );
  XOR2_X1 U759 ( .A(n458), .B(KEYINPUT127), .Z(n712) );
  XNOR2_X1 U760 ( .A(n711), .B(n712), .ZN(n716) );
  XNOR2_X1 U761 ( .A(n713), .B(n716), .ZN(n715) );
  NAND2_X1 U762 ( .A1(n715), .A2(n714), .ZN(n720) );
  XNOR2_X1 U763 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(G900), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n718), .A2(G953), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n720), .A2(n719), .ZN(G72) );
  XOR2_X1 U767 ( .A(G122), .B(n721), .Z(G24) );
  XOR2_X1 U768 ( .A(G137), .B(n722), .Z(G39) );
  XNOR2_X1 U769 ( .A(G119), .B(n723), .ZN(G21) );
  XOR2_X1 U770 ( .A(n724), .B(G131), .Z(G33) );
endmodule

