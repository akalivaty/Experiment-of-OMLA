//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT28), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n216), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n218), .A2(new_n214), .A3(new_n215), .A4(KEYINPUT67), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n217), .A2(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n213), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT68), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n214), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT25), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(G183gat), .B(G190gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n233), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT66), .B(G169gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n230), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n229), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(new_n236), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n222), .A2(new_n226), .B1(new_n237), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n202), .B1(new_n243), .B2(KEYINPUT29), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G197gat), .B(G204gat), .Z(new_n247));
  AND2_X1   g046(.A1(G211gat), .A2(G218gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(KEYINPUT22), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n247), .B2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n242), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n220), .A2(new_n221), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n221), .A3(new_n224), .ZN(new_n257));
  INV_X1    g056(.A(new_n213), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n255), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n202), .B(KEYINPUT78), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(KEYINPUT79), .B(new_n202), .C1(new_n243), .C2(KEYINPUT29), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n246), .A2(new_n254), .A3(new_n262), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n254), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT29), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n243), .A2(new_n202), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT80), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n273), .A3(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT30), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n264), .A2(new_n282), .A3(new_n273), .A4(new_n269), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G127gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G134gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G127gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g090(.A1(G113gat), .A2(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G113gat), .A2(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G113gat), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n292), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n290), .A2(new_n295), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G141gat), .B(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n307), .B(new_n306), .C1(new_n302), .C2(KEYINPUT2), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n287), .B2(new_n289), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n288), .A2(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n286), .A2(G134gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n293), .B2(new_n294), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n298), .A2(KEYINPUT70), .A3(new_n292), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n300), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n319), .A2(new_n323), .A3(KEYINPUT71), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT71), .B1(new_n319), .B2(new_n323), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n301), .B(new_n313), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n301), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n323), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n323), .A3(KEYINPUT71), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n312), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n311), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n326), .B(KEYINPUT4), .C1(new_n332), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT39), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n332), .A2(new_n341), .A3(new_n313), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n338), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT0), .ZN(new_n345));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  AND2_X1   g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  OR3_X1    g147(.A1(new_n332), .A2(KEYINPUT82), .A3(new_n313), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n301), .B1(new_n324), .B2(new_n325), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n312), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n326), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n342), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT39), .B1(new_n354), .B2(new_n339), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT40), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n347), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n349), .A2(new_n352), .A3(KEYINPUT5), .A4(new_n340), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT81), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n354), .B2(new_n339), .ZN(new_n364));
  AOI211_X1 g163(.A(new_n340), .B(new_n362), .C1(new_n337), .C2(new_n342), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n359), .B(new_n360), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n356), .B2(new_n357), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n285), .A2(new_n358), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n280), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n264), .A2(new_n269), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n274), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT37), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n267), .A2(new_n268), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n254), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n246), .A2(new_n265), .A3(new_n262), .A4(new_n263), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT38), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n370), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OR3_X1    g181(.A1(new_n381), .A2(new_n382), .A3(new_n347), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n264), .B2(new_n269), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT38), .B1(new_n373), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n347), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n382), .A3(new_n366), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n380), .A2(new_n383), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT31), .B(G50gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n252), .B2(new_n253), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n312), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT85), .ZN(new_n395));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n335), .A2(new_n266), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n265), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n312), .C1(new_n393), .C2(KEYINPUT3), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n395), .A2(new_n397), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n253), .A2(KEYINPUT83), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT29), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n252), .A2(KEYINPUT83), .A3(new_n253), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(KEYINPUT84), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n334), .A3(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n410), .A2(new_n312), .B1(new_n265), .B2(new_n398), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n411), .B2(new_n397), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(G22gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n392), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n402), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n409), .A2(new_n334), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT84), .B1(new_n404), .B2(new_n405), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n312), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n399), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n416), .B1(new_n420), .B2(new_n396), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(G22gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n391), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n412), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n369), .A2(new_n388), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT36), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT34), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(KEYINPUT64), .Z(new_n434));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n350), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(KEYINPUT73), .B(new_n301), .C1(new_n324), .C2(new_n325), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n260), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n243), .A2(new_n435), .A3(new_n350), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(KEYINPUT76), .A3(new_n439), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n432), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n434), .B(KEYINPUT65), .Z(new_n445));
  AOI211_X1 g244(.A(KEYINPUT34), .B(new_n445), .C1(new_n438), .C2(new_n439), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT77), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  INV_X1    g248(.A(new_n443), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT76), .B1(new_n438), .B2(new_n439), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(new_n451), .A3(new_n434), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n448), .B(new_n449), .C1(new_n452), .C2(new_n432), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n439), .A3(new_n445), .ZN(new_n454));
  XOR2_X1   g253(.A(G15gat), .B(G43gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT74), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT33), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n454), .A2(KEYINPUT75), .A3(KEYINPUT32), .A4(new_n459), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n458), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n454), .B2(KEYINPUT32), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n462), .A2(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n447), .A2(new_n453), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n447), .B2(new_n453), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n431), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n440), .A2(new_n441), .ZN(new_n473));
  INV_X1    g272(.A(new_n434), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n443), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT34), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n448), .B1(new_n476), .B2(new_n449), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n444), .A2(KEYINPUT77), .A3(new_n446), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n447), .A2(new_n453), .A3(new_n468), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT36), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n423), .A2(new_n415), .B1(new_n426), .B2(new_n427), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n387), .A2(new_n383), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n276), .A2(new_n278), .B1(new_n281), .B2(new_n283), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n471), .A2(new_n481), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n469), .A2(new_n470), .A3(new_n482), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n483), .A2(KEYINPUT89), .A3(new_n484), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n429), .A3(new_n480), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT89), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n430), .A2(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G57gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT95), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G57gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n498), .A3(G64gat), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n495), .A2(G64gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT96), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(KEYINPUT96), .A3(new_n500), .ZN(new_n504));
  INV_X1    g303(.A(G71gat), .ZN(new_n505));
  INV_X1    g304(.A(G78gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT9), .ZN(new_n508));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512));
  OAI22_X1  g311(.A1(new_n512), .A2(KEYINPUT94), .B1(KEYINPUT9), .B2(new_n507), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n512), .A2(KEYINPUT94), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT98), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(KEYINPUT21), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n522), .A3(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G8gat), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(new_n531), .A3(new_n526), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n520), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT21), .B1(new_n511), .B2(new_n515), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  XNOR2_X1  g341(.A(G127gat), .B(G155gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT20), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n542), .A2(new_n544), .ZN(new_n547));
  XOR2_X1   g346(.A(G183gat), .B(G211gat), .Z(new_n548));
  NOR3_X1   g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n542), .A2(new_n544), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n539), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n546), .B2(new_n547), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n550), .A3(new_n545), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n537), .A4(new_n538), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G92gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT100), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G99gat), .A3(G106gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n569), .A3(new_n571), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n564), .A2(new_n571), .A3(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT101), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  OR2_X1    g382(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n585));
  AOI21_X1  g384(.A(G36gat), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G29gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT15), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G43gat), .B(G50gat), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT15), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n584), .A2(new_n585), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n593), .B(new_n588), .C1(new_n594), .C2(G36gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n590), .A3(new_n591), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n583), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n592), .A2(new_n596), .A3(new_n583), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n582), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n571), .B1(new_n564), .B2(new_n569), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n578), .A2(new_n602), .A3(KEYINPUT101), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n575), .A2(new_n574), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT102), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n596), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n599), .A2(new_n601), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n612), .A2(KEYINPUT103), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n599), .A2(new_n609), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n600), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(KEYINPUT103), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G134gat), .B(G162gat), .Z(new_n618));
  NOR2_X1   g417(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n614), .B2(new_n600), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n617), .A2(new_n621), .B1(new_n612), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n558), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n511), .A2(new_n518), .A3(new_n515), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n518), .B1(new_n511), .B2(new_n515), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n607), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n576), .A2(new_n579), .B1(new_n511), .B2(new_n515), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n573), .A2(new_n575), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n633), .A2(new_n515), .A3(new_n511), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n629), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI211_X1 g434(.A(KEYINPUT104), .B(new_n626), .C1(new_n631), .C2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n517), .A2(KEYINPUT10), .A3(new_n519), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n582), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n639), .B2(new_n625), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n516), .B1(new_n603), .B2(new_n604), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n633), .A2(new_n511), .A3(new_n515), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n626), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT105), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n646), .A2(new_n650), .A3(new_n626), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT106), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n645), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n626), .B1(new_n631), .B2(new_n635), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n645), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n661));
  NAND2_X1  g460(.A1(G229gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AND4_X1   g462(.A1(new_n530), .A2(new_n532), .A3(new_n596), .A4(new_n592), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n530), .A2(new_n532), .B1(new_n592), .B2(new_n596), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT93), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT93), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n668), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n534), .B1(new_n598), .B2(new_n597), .ZN(new_n671));
  INV_X1    g470(.A(new_n665), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n662), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n671), .A2(KEYINPUT18), .A3(new_n672), .A4(new_n662), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(G169gat), .B(G197gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT12), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n670), .A2(new_n675), .A3(new_n676), .A4(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OR4_X1    g487(.A1(new_n494), .A2(new_n624), .A3(new_n660), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n483), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n524), .ZN(G1324gat));
  NOR2_X1   g490(.A1(new_n689), .A2(new_n484), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n531), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT16), .B(G8gat), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n689), .A2(new_n484), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n471), .A2(new_n481), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n689), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n469), .A2(new_n470), .ZN(new_n700));
  INV_X1    g499(.A(G15gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n689), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n429), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n494), .B2(new_n623), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n490), .A2(new_n493), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n485), .A2(new_n482), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n698), .A2(new_n430), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n623), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(KEYINPUT44), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n558), .A2(new_n660), .A3(new_n688), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n483), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n623), .B1(new_n710), .B2(new_n712), .ZN(new_n720));
  INV_X1    g519(.A(new_n483), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n720), .A2(new_n587), .A3(new_n721), .A4(new_n717), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT108), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n719), .B1(new_n724), .B2(new_n725), .ZN(G1328gat));
  NAND2_X1  g525(.A1(new_n720), .A2(new_n717), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(G36gat), .A3(new_n484), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT46), .ZN(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n718), .B2(new_n484), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n698), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n709), .A2(new_n715), .A3(new_n732), .A4(new_n717), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n735), .A3(new_n700), .A4(new_n717), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n737), .B(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n720), .A2(KEYINPUT110), .A3(new_n717), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n429), .A2(G50gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n709), .A2(new_n715), .A3(new_n482), .A4(new_n717), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT112), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(KEYINPUT112), .ZN(new_n749));
  OAI211_X1 g548(.A(KEYINPUT48), .B(new_n745), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(G50gat), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT48), .B1(new_n751), .B2(new_n745), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n754), .B(KEYINPUT48), .C1(new_n751), .C2(new_n745), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n753), .B2(new_n755), .ZN(G1331gat));
  INV_X1    g555(.A(new_n660), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n624), .A2(new_n757), .A3(new_n687), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n713), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n721), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n496), .A2(new_n498), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1332gat));
  NOR2_X1   g562(.A1(new_n759), .A2(new_n484), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n765), .ZN(G1333gat));
  OAI21_X1  g567(.A(G71gat), .B1(new_n759), .B2(new_n698), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n700), .A2(new_n505), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g571(.A1(new_n759), .A2(new_n429), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n506), .ZN(G1335gat));
  NOR3_X1   g573(.A1(new_n558), .A2(new_n757), .A3(new_n687), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n716), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n483), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n558), .A2(new_n687), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n720), .B2(new_n778), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n483), .A2(new_n757), .A3(G85gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(G1336gat));
  NAND4_X1  g583(.A1(new_n709), .A2(new_n715), .A3(new_n285), .A4(new_n775), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n285), .A2(new_n559), .A3(new_n660), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT113), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n779), .B2(new_n780), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n776), .B2(new_n698), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n757), .A2(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n781), .A2(new_n700), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n709), .A2(new_n715), .A3(new_n482), .A4(new_n775), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n757), .A2(new_n429), .A3(G106gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n779), .B2(new_n780), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n796), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT115), .B(new_n800), .C1(new_n779), .C2(new_n780), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n809), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n808), .B(new_n801), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n807), .A2(new_n813), .ZN(G1339gat));
  NOR2_X1   g613(.A1(new_n285), .A2(new_n483), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n635), .B(new_n626), .C1(new_n582), .C2(new_n638), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n636), .A2(new_n640), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n639), .A2(new_n625), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT55), .B(new_n645), .C1(new_n821), .C2(KEYINPUT54), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(KEYINPUT104), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n639), .A2(new_n637), .A3(new_n625), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n649), .A2(new_n654), .A3(new_n651), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n654), .B1(new_n649), .B2(new_n651), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n644), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n820), .A2(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n646), .A2(new_n647), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n630), .A2(new_n607), .B1(new_n831), .B2(new_n629), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n832), .B2(new_n626), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n823), .A2(new_n833), .A3(new_n824), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n644), .B1(new_n658), .B2(new_n830), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n817), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n838), .B(new_n644), .C1(new_n658), .C2(new_n830), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n834), .A2(new_n839), .B1(new_n641), .B2(new_n656), .ZN(new_n840));
  INV_X1    g639(.A(new_n835), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n820), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT118), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n843), .A3(new_n687), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n662), .B1(new_n671), .B2(new_n672), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n664), .A2(new_n665), .A3(new_n663), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n682), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n686), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n657), .B2(new_n659), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n714), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n848), .B(KEYINPUT119), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n714), .A2(new_n837), .A3(new_n843), .A4(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n557), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n558), .A2(new_n623), .A3(new_n757), .A4(new_n688), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n816), .B1(new_n858), .B2(new_n429), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT120), .B(new_n482), .C1(new_n854), .C2(new_n857), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n700), .B(new_n815), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n296), .A3(new_n688), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n483), .B1(new_n854), .B2(new_n857), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(new_n484), .A3(new_n487), .ZN(new_n864));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n687), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n297), .A3(new_n660), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n859), .A2(new_n860), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n700), .A3(new_n660), .A4(new_n815), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT121), .B1(new_n869), .B2(G120gat), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT121), .B(G120gat), .C1(new_n861), .C2(new_n757), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n861), .B2(new_n557), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n864), .A2(new_n286), .A3(new_n558), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1342gat));
  OAI21_X1  g675(.A(G134gat), .B1(new_n861), .B2(new_n623), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n623), .A2(new_n285), .A3(G134gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n487), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT122), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n877), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n698), .A2(new_n815), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n858), .B2(new_n482), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n842), .A2(KEYINPUT123), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n836), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n893), .A3(new_n687), .A4(new_n840), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n714), .B1(new_n894), .B2(new_n850), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n557), .B1(new_n895), .B2(new_n853), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n890), .B(new_n429), .C1(new_n896), .C2(new_n857), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n888), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G141gat), .B1(new_n898), .B2(new_n688), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n863), .A2(new_n482), .A3(new_n698), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n484), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n688), .A2(G141gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n899), .B(new_n905), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n898), .A2(new_n757), .ZN(new_n908));
  INV_X1    g707(.A(G148gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n660), .B1(new_n888), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n912), .B2(new_n888), .ZN(new_n914));
  INV_X1    g713(.A(new_n855), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n714), .A2(new_n852), .A3(new_n840), .A4(new_n842), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n839), .A2(new_n834), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n687), .A3(new_n657), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT123), .B(KEYINPUT55), .C1(new_n834), .C2(new_n835), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n849), .B1(new_n920), .B2(new_n891), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n916), .B1(new_n921), .B2(new_n714), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(new_n557), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n890), .B1(new_n923), .B2(new_n429), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n429), .B1(new_n854), .B2(new_n857), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n924), .A2(new_n925), .B1(KEYINPUT57), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n925), .A3(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n914), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n911), .B1(new_n930), .B2(G148gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n660), .A2(new_n909), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n910), .A2(new_n931), .B1(new_n901), .B2(new_n932), .ZN(G1345gat));
  OAI21_X1  g732(.A(G155gat), .B1(new_n898), .B2(new_n557), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n558), .A2(new_n304), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n901), .B2(new_n935), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n898), .B2(new_n623), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n900), .A2(new_n305), .A3(new_n484), .A4(new_n714), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n721), .A2(new_n484), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n700), .B(new_n940), .C1(new_n859), .C2(new_n860), .ZN(new_n941));
  OAI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n688), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n721), .B1(new_n854), .B2(new_n857), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(new_n285), .A3(new_n487), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n239), .A3(new_n687), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1348gat));
  OAI21_X1  g749(.A(G176gat), .B1(new_n941), .B2(new_n757), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n944), .A2(new_n215), .A3(new_n660), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1349gat));
  OAI21_X1  g752(.A(G183gat), .B1(new_n941), .B2(new_n557), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n210), .A3(new_n558), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT127), .B(KEYINPUT60), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n207), .A3(new_n714), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n868), .A2(new_n700), .A3(new_n714), .A4(new_n940), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(G190gat), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n963), .B(G190gat), .C1(new_n941), .C2(new_n623), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n962), .B1(new_n965), .B2(new_n967), .ZN(G1351gat));
  NOR3_X1   g767(.A1(new_n732), .A2(new_n429), .A3(new_n484), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n943), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n687), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n698), .A2(new_n940), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n924), .A2(new_n925), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n926), .A2(KEYINPUT57), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n976), .B2(new_n928), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n687), .A2(G197gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(G1352gat));
  NOR3_X1   g778(.A1(new_n970), .A2(G204gat), .A3(new_n757), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT62), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n977), .A2(new_n660), .ZN(new_n982));
  INV_X1    g781(.A(G204gat), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(G1353gat));
  OR3_X1    g783(.A1(new_n970), .A2(G211gat), .A3(new_n557), .ZN(new_n985));
  INV_X1    g784(.A(new_n973), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n558), .B(new_n986), .C1(new_n927), .C2(new_n929), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  INV_X1    g789(.A(G218gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n991), .A3(new_n714), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n977), .A2(new_n714), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(new_n991), .ZN(G1355gat));
endmodule


