

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n722), .A2(n721), .ZN(n748) );
  XOR2_X2 U555 ( .A(KEYINPUT64), .B(n527), .Z(n903) );
  XNOR2_X1 U556 ( .A(n755), .B(n754), .ZN(n785) );
  INV_X2 U557 ( .A(n748), .ZN(n767) );
  INV_X1 U558 ( .A(n720), .ZN(n721) );
  NOR2_X1 U559 ( .A1(n786), .A2(n785), .ZN(n522) );
  INV_X1 U560 ( .A(G8), .ZN(n756) );
  NOR2_X1 U561 ( .A1(n778), .A2(n756), .ZN(n757) );
  INV_X1 U562 ( .A(KEYINPUT103), .ZN(n796) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  AND2_X1 U564 ( .A1(n813), .A2(n812), .ZN(n815) );
  NOR2_X1 U565 ( .A1(G651), .A2(n648), .ZN(n642) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n632) );
  XNOR2_X1 U567 ( .A(n532), .B(KEYINPUT92), .ZN(G164) );
  INV_X1 U568 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n526), .ZN(n901) );
  NAND2_X1 U570 ( .A1(G126), .A2(n901), .ZN(n525) );
  XOR2_X2 U571 ( .A(KEYINPUT17), .B(n523), .Z(n898) );
  NAND2_X1 U572 ( .A1(G138), .A2(n898), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n531) );
  AND2_X1 U574 ( .A1(n526), .A2(G2104), .ZN(n897) );
  NAND2_X1 U575 ( .A1(G102), .A2(n897), .ZN(n529) );
  NAND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  NAND2_X1 U577 ( .A1(G114), .A2(n903), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U580 ( .A(G651), .ZN(n538) );
  NOR2_X1 U581 ( .A1(G543), .A2(n538), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n533), .Z(n646) );
  NAND2_X1 U583 ( .A1(G63), .A2(n646), .ZN(n535) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  NAND2_X1 U585 ( .A1(G51), .A2(n642), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U587 ( .A(KEYINPUT6), .B(n536), .ZN(n544) );
  NAND2_X1 U588 ( .A1(n632), .A2(G89), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n537), .B(KEYINPUT4), .ZN(n540) );
  NOR2_X1 U590 ( .A1(n648), .A2(n538), .ZN(n635) );
  NAND2_X1 U591 ( .A1(G76), .A2(n635), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U593 ( .A(KEYINPUT75), .B(n541), .ZN(n542) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n542), .ZN(n543) );
  NOR2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n545), .Z(G168) );
  XOR2_X1 U597 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U598 ( .A1(G75), .A2(n635), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G88), .A2(n632), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n552) );
  NAND2_X1 U601 ( .A1(G62), .A2(n646), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G50), .A2(n642), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U604 ( .A(KEYINPUT83), .B(n550), .Z(n551) );
  NOR2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U606 ( .A(KEYINPUT84), .B(n553), .ZN(G166) );
  INV_X1 U607 ( .A(G166), .ZN(G303) );
  NAND2_X1 U608 ( .A1(G64), .A2(n646), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G52), .A2(n642), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n562) );
  NAND2_X1 U611 ( .A1(n635), .A2(G77), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT66), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G90), .A2(n632), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(KEYINPUT9), .B(n559), .ZN(n560) );
  XNOR2_X1 U616 ( .A(KEYINPUT67), .B(n560), .ZN(n561) );
  NOR2_X1 U617 ( .A1(n562), .A2(n561), .ZN(G171) );
  INV_X1 U618 ( .A(G171), .ZN(G301) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U620 ( .A(G69), .ZN(G235) );
  INV_X1 U621 ( .A(G108), .ZN(G238) );
  INV_X1 U622 ( .A(G120), .ZN(G236) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n563) );
  XOR2_X1 U626 ( .A(n563), .B(KEYINPUT10), .Z(n833) );
  AND2_X1 U627 ( .A1(G567), .A2(n833), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT11), .ZN(G234) );
  XNOR2_X1 U629 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n635), .A2(G68), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT71), .B(n566), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n632), .A2(G81), .ZN(n567) );
  XOR2_X1 U634 ( .A(n567), .B(KEYINPUT12), .Z(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(n574) );
  NAND2_X1 U637 ( .A1(n646), .A2(G56), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n642), .A2(G43), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n734) );
  INV_X1 U642 ( .A(n734), .ZN(n929) );
  NAND2_X1 U643 ( .A1(n929), .A2(G860), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G79), .A2(n635), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G92), .A2(n632), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G66), .A2(n646), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G54), .A2(n642), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n583), .Z(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT74), .B(n584), .Z(n602) );
  NOR2_X1 U653 ( .A1(n602), .A2(G868), .ZN(n586) );
  INV_X1 U654 ( .A(G868), .ZN(n663) );
  NOR2_X1 U655 ( .A1(n663), .A2(G301), .ZN(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G78), .A2(n635), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT68), .B(n587), .Z(n592) );
  NAND2_X1 U659 ( .A1(G65), .A2(n646), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G53), .A2(n642), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT69), .B(n590), .Z(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n632), .A2(G91), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(G299) );
  XOR2_X1 U666 ( .A(KEYINPUT76), .B(G868), .Z(n595) );
  NOR2_X1 U667 ( .A1(G286), .A2(n595), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT77), .B(n596), .Z(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U671 ( .A(KEYINPUT78), .B(n599), .ZN(G297) );
  INV_X1 U672 ( .A(G559), .ZN(n600) );
  NOR2_X1 U673 ( .A1(G860), .A2(n600), .ZN(n601) );
  XNOR2_X1 U674 ( .A(KEYINPUT79), .B(n601), .ZN(n603) );
  INV_X1 U675 ( .A(n602), .ZN(n937) );
  NAND2_X1 U676 ( .A1(n603), .A2(n937), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n734), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n937), .A2(G868), .ZN(n605) );
  NOR2_X1 U680 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U681 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n897), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G111), .A2(n903), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U685 ( .A(KEYINPUT80), .B(n610), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n901), .A2(G123), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G135), .A2(n898), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n1002) );
  XNOR2_X1 U691 ( .A(G2096), .B(n1002), .ZN(n616) );
  INV_X1 U692 ( .A(G2100), .ZN(n870) );
  NAND2_X1 U693 ( .A1(n616), .A2(n870), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n937), .ZN(n660) );
  XOR2_X1 U695 ( .A(n929), .B(n660), .Z(n617) );
  NOR2_X1 U696 ( .A1(n617), .A2(G860), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G80), .A2(n635), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G93), .A2(n632), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G67), .A2(n646), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G55), .A2(n642), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n662) );
  XOR2_X1 U704 ( .A(n624), .B(n662), .Z(G145) );
  NAND2_X1 U705 ( .A1(G60), .A2(n646), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G47), .A2(n642), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U708 ( .A(KEYINPUT65), .B(n627), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G72), .A2(n635), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G85), .A2(n632), .ZN(n628) );
  AND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G86), .A2(n632), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G61), .A2(n646), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G48), .A2(n642), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n642), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT81), .B(n647), .Z(n650) );
  NAND2_X1 U727 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(G288) );
  XOR2_X1 U729 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n652) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n652), .B(n651), .ZN(n656) );
  XOR2_X1 U732 ( .A(G299), .B(G303), .Z(n654) );
  XNOR2_X1 U733 ( .A(G290), .B(G305), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(n658) );
  XOR2_X1 U736 ( .A(G288), .B(n662), .Z(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U738 ( .A(n659), .B(n929), .Z(n919) );
  XNOR2_X1 U739 ( .A(n660), .B(n919), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U749 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U752 ( .A1(G218), .A2(n671), .ZN(n672) );
  XNOR2_X1 U753 ( .A(KEYINPUT88), .B(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G96), .ZN(n674) );
  XOR2_X1 U755 ( .A(KEYINPUT89), .B(n674), .Z(n838) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n838), .ZN(n675) );
  XOR2_X1 U757 ( .A(KEYINPUT90), .B(n675), .Z(n680) );
  NOR2_X1 U758 ( .A1(G236), .A2(G238), .ZN(n677) );
  NOR2_X1 U759 ( .A1(G235), .A2(G237), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U761 ( .A(KEYINPUT91), .B(n678), .Z(n839) );
  AND2_X1 U762 ( .A1(n839), .A2(G567), .ZN(n679) );
  NOR2_X1 U763 ( .A1(n680), .A2(n679), .ZN(G319) );
  INV_X1 U764 ( .A(G319), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n837) );
  NAND2_X1 U767 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U768 ( .A1(G113), .A2(n903), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G101), .A2(n897), .ZN(n683) );
  XOR2_X1 U770 ( .A(KEYINPUT23), .B(n683), .Z(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U772 ( .A1(G125), .A2(n901), .ZN(n687) );
  NAND2_X1 U773 ( .A1(G137), .A2(n898), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U775 ( .A1(n689), .A2(n688), .ZN(G160) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n722), .A2(n720), .ZN(n827) );
  INV_X1 U779 ( .A(G2067), .ZN(n867) );
  XOR2_X1 U780 ( .A(n867), .B(KEYINPUT37), .Z(n816) );
  NAND2_X1 U781 ( .A1(G104), .A2(n897), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G140), .A2(n898), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U784 ( .A(KEYINPUT34), .B(n692), .ZN(n698) );
  NAND2_X1 U785 ( .A1(G116), .A2(n903), .ZN(n693) );
  XOR2_X1 U786 ( .A(KEYINPUT93), .B(n693), .Z(n695) );
  NAND2_X1 U787 ( .A1(n901), .A2(G128), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U789 ( .A(KEYINPUT35), .B(n696), .Z(n697) );
  NOR2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U791 ( .A(KEYINPUT36), .B(n699), .ZN(n909) );
  NOR2_X1 U792 ( .A1(n816), .A2(n909), .ZN(n1017) );
  NAND2_X1 U793 ( .A1(n827), .A2(n1017), .ZN(n824) );
  NAND2_X1 U794 ( .A1(n901), .A2(G119), .ZN(n701) );
  NAND2_X1 U795 ( .A1(G107), .A2(n903), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n897), .A2(G95), .ZN(n702) );
  XOR2_X1 U798 ( .A(KEYINPUT94), .B(n702), .Z(n703) );
  NOR2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n898), .A2(G131), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n912) );
  AND2_X1 U802 ( .A1(n912), .A2(G1991), .ZN(n717) );
  NAND2_X1 U803 ( .A1(G141), .A2(n898), .ZN(n707) );
  XNOR2_X1 U804 ( .A(n707), .B(KEYINPUT96), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n897), .A2(G105), .ZN(n708) );
  XNOR2_X1 U806 ( .A(n708), .B(KEYINPUT38), .ZN(n710) );
  NAND2_X1 U807 ( .A1(G129), .A2(n901), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U809 ( .A1(G117), .A2(n903), .ZN(n711) );
  XNOR2_X1 U810 ( .A(KEYINPUT95), .B(n711), .ZN(n712) );
  NOR2_X1 U811 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n913) );
  AND2_X1 U813 ( .A1(n913), .A2(G1996), .ZN(n716) );
  NOR2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n1008) );
  INV_X1 U815 ( .A(n1008), .ZN(n718) );
  NAND2_X1 U816 ( .A1(n718), .A2(n827), .ZN(n817) );
  NAND2_X1 U817 ( .A1(n824), .A2(n817), .ZN(n719) );
  XNOR2_X1 U818 ( .A(KEYINPUT97), .B(n719), .ZN(n813) );
  INV_X1 U819 ( .A(G299), .ZN(n729) );
  NAND2_X1 U820 ( .A1(G1956), .A2(n767), .ZN(n723) );
  XNOR2_X1 U821 ( .A(KEYINPUT99), .B(n723), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n748), .A2(G2072), .ZN(n724) );
  XNOR2_X1 U823 ( .A(KEYINPUT27), .B(n724), .ZN(n725) );
  NOR2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n727) );
  XOR2_X1 U826 ( .A(n727), .B(KEYINPUT28), .Z(n746) );
  NAND2_X1 U827 ( .A1(n729), .A2(n728), .ZN(n744) );
  AND2_X1 U828 ( .A1(n748), .A2(G1996), .ZN(n730) );
  XOR2_X1 U829 ( .A(n730), .B(KEYINPUT26), .Z(n732) );
  NAND2_X1 U830 ( .A1(n767), .A2(G1341), .ZN(n731) );
  NAND2_X1 U831 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U832 ( .A1(n734), .A2(n733), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n937), .A2(n740), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n767), .A2(n867), .ZN(n735) );
  XOR2_X1 U835 ( .A(n735), .B(KEYINPUT100), .Z(n737) );
  NAND2_X1 U836 ( .A1(n767), .A2(G1348), .ZN(n736) );
  NAND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U838 ( .A1(n739), .A2(n738), .ZN(n742) );
  OR2_X1 U839 ( .A1(n937), .A2(n740), .ZN(n741) );
  NAND2_X1 U840 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U843 ( .A(n747), .B(KEYINPUT29), .ZN(n752) );
  NAND2_X1 U844 ( .A1(G1961), .A2(n767), .ZN(n750) );
  XOR2_X1 U845 ( .A(KEYINPUT25), .B(G2078), .Z(n960) );
  NAND2_X1 U846 ( .A1(n748), .A2(n960), .ZN(n749) );
  NAND2_X1 U847 ( .A1(n750), .A2(n749), .ZN(n753) );
  NOR2_X1 U848 ( .A1(G301), .A2(n753), .ZN(n751) );
  NOR2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n765) );
  AND2_X1 U850 ( .A1(G301), .A2(n753), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n767), .A2(G8), .ZN(n755) );
  INV_X1 U852 ( .A(KEYINPUT98), .ZN(n754) );
  INV_X1 U853 ( .A(n785), .ZN(n807) );
  NOR2_X2 U854 ( .A1(n807), .A2(G1966), .ZN(n777) );
  INV_X1 U855 ( .A(n777), .ZN(n758) );
  NOR2_X1 U856 ( .A1(G2084), .A2(n767), .ZN(n778) );
  NAND2_X1 U857 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U858 ( .A(KEYINPUT30), .B(n759), .ZN(n760) );
  NOR2_X1 U859 ( .A1(G168), .A2(n760), .ZN(n761) );
  NOR2_X1 U860 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U861 ( .A(n763), .B(KEYINPUT31), .ZN(n764) );
  NOR2_X1 U862 ( .A1(n765), .A2(n764), .ZN(n776) );
  INV_X1 U863 ( .A(n776), .ZN(n766) );
  NAND2_X1 U864 ( .A1(n766), .A2(G286), .ZN(n773) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n767), .ZN(n768) );
  XNOR2_X1 U866 ( .A(n768), .B(KEYINPUT102), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n807), .A2(G1971), .ZN(n769) );
  NOR2_X1 U868 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n771), .A2(G303), .ZN(n772) );
  NAND2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U871 ( .A1(n774), .A2(G8), .ZN(n775) );
  XNOR2_X1 U872 ( .A(n775), .B(KEYINPUT32), .ZN(n800) );
  NOR2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U874 ( .A1(G8), .A2(n778), .ZN(n779) );
  AND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U876 ( .A(n781), .B(KEYINPUT101), .ZN(n799) );
  INV_X1 U877 ( .A(KEYINPUT33), .ZN(n782) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n936) );
  AND2_X1 U879 ( .A1(n782), .A2(n936), .ZN(n787) );
  AND2_X1 U880 ( .A1(n799), .A2(n787), .ZN(n783) );
  NAND2_X1 U881 ( .A1(n800), .A2(n783), .ZN(n795) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n789), .A2(n785), .ZN(n784) );
  NAND2_X1 U884 ( .A1(n784), .A2(KEYINPUT33), .ZN(n791) );
  INV_X1 U885 ( .A(n791), .ZN(n786) );
  INV_X1 U886 ( .A(n787), .ZN(n790) );
  NOR2_X1 U887 ( .A1(G303), .A2(G1971), .ZN(n788) );
  NOR2_X1 U888 ( .A1(n789), .A2(n788), .ZN(n931) );
  OR2_X1 U889 ( .A1(n790), .A2(n931), .ZN(n792) );
  AND2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  OR2_X1 U891 ( .A1(n522), .A2(n793), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n797) );
  XNOR2_X1 U893 ( .A(n797), .B(n796), .ZN(n798) );
  XOR2_X1 U894 ( .A(G1981), .B(G305), .Z(n932) );
  NAND2_X1 U895 ( .A1(n798), .A2(n932), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n803) );
  NOR2_X1 U897 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U898 ( .A1(G8), .A2(n801), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U900 ( .A1(n807), .A2(n804), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XOR2_X1 U902 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n947) );
  NAND2_X1 U907 ( .A1(n947), .A2(n827), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n830) );
  NAND2_X1 U909 ( .A1(n816), .A2(n909), .ZN(n1014) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n913), .ZN(n1010) );
  INV_X1 U911 ( .A(n817), .ZN(n820) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n912), .ZN(n1003) );
  NOR2_X1 U914 ( .A1(n818), .A2(n1003), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n1010), .A2(n821), .ZN(n822) );
  XNOR2_X1 U917 ( .A(KEYINPUT39), .B(n822), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT104), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n1014), .A2(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U924 ( .A1(n833), .A2(G2106), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT109), .B(n832), .Z(G217) );
  INV_X1 U926 ( .A(n833), .ZN(G223) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT110), .B(n834), .Z(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U932 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT105), .B(KEYINPUT107), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2446), .B(G2451), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(n842), .B(G2430), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT106), .B(G2438), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2435), .B(G2454), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2443), .B(G2427), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G14), .A2(n851), .ZN(n852) );
  XOR2_X1 U949 ( .A(KEYINPUT108), .B(n852), .Z(G401) );
  XOR2_X1 U950 ( .A(G2474), .B(G1986), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(KEYINPUT113), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1976), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(G1956), .B(G1961), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1981), .B(G1966), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G229) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT112), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2090), .B(KEYINPUT43), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U965 ( .A(n866), .B(KEYINPUT42), .Z(n869) );
  XOR2_X1 U966 ( .A(n867), .B(G2072), .Z(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n874) );
  XNOR2_X1 U968 ( .A(G2678), .B(n870), .ZN(n872) );
  XNOR2_X1 U969 ( .A(G2078), .B(G2084), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(G227) );
  NAND2_X1 U972 ( .A1(G124), .A2(n901), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT115), .B(n875), .Z(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G100), .A2(n897), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U977 ( .A1(n898), .A2(G136), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G112), .A2(n903), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(KEYINPUT116), .B(n883), .ZN(G162) );
  NAND2_X1 U982 ( .A1(n901), .A2(G130), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G118), .A2(n903), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n892) );
  XNOR2_X1 U985 ( .A(KEYINPUT118), .B(KEYINPUT45), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n898), .A2(G142), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n897), .A2(G106), .ZN(n886) );
  XOR2_X1 U988 ( .A(KEYINPUT117), .B(n886), .Z(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n894) );
  XNOR2_X1 U993 ( .A(G160), .B(n1002), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n911) );
  NAND2_X1 U996 ( .A1(G103), .A2(n897), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G139), .A2(n898), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n908) );
  NAND2_X1 U999 ( .A1(n901), .A2(G127), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT119), .B(n902), .Z(n905) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n903), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n906), .Z(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n998) );
  XNOR2_X1 U1005 ( .A(n909), .B(n998), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n917) );
  XOR2_X1 U1007 ( .A(n913), .B(n912), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(G162), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(G164), .B(n915), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1012 ( .A(n937), .B(G286), .Z(n920) );
  XNOR2_X1 U1013 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1014 ( .A(n921), .B(G301), .Z(n922) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n922), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G229), .A2(G227), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n924), .ZN(n925) );
  AND2_X1 U1019 ( .A1(G319), .A2(n925), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1023 ( .A(KEYINPUT56), .B(G16), .ZN(n951) );
  XOR2_X1 U1024 ( .A(G1341), .B(KEYINPUT124), .Z(n928) );
  XOR2_X1 U1025 ( .A(n929), .B(n928), .Z(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n943) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(n934), .B(KEYINPUT57), .ZN(n941) );
  NAND2_X1 U1030 ( .A1(G303), .A2(G1971), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1032 ( .A(G1348), .B(n937), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G299), .B(G1956), .Z(n945) );
  XOR2_X1 U1037 ( .A(G301), .B(G1961), .Z(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n1030) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n959) );
  XOR2_X1 U1045 ( .A(G26), .B(G2067), .Z(n954) );
  NAND2_X1 U1046 ( .A1(n954), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G25), .B(G1991), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT122), .B(n955), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G27), .B(n960), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(KEYINPUT123), .B(n963), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n964), .B(KEYINPUT53), .ZN(n969) );
  XNOR2_X1 U1055 ( .A(G2084), .B(G34), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n965), .B(KEYINPUT54), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n970), .Z(n972) );
  INV_X1 U1061 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n973), .ZN(n1028) );
  XOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .Z(n974) );
  XNOR2_X1 U1065 ( .A(G4), .B(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G20), .B(G1956), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(KEYINPUT60), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G24), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G22), .B(G1971), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G1976), .B(KEYINPUT125), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n984), .B(G23), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G21), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G1961), .B(G5), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(KEYINPUT61), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT126), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(G16), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(KEYINPUT127), .B(n997), .ZN(n1026) );
  XOR2_X1 U1089 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1001), .Z(n1020) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1004), .Z(n1006) );
  XOR2_X1 U1095 ( .A(G2084), .B(G160), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT51), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT121), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1031), .ZN(G150) );
  INV_X1 U1114 ( .A(G150), .ZN(G311) );
endmodule

