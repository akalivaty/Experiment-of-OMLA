//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT64), .Z(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n210), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n219), .B1(new_n213), .B2(new_n212), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT67), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n214), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(new_n257), .B2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G223), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n261), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G222), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n258), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G200), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n215), .A2(G33), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n214), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n281), .A2(new_n286), .B1(new_n202), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n250), .B2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT9), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n276), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT73), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  OAI211_X1 g0096(.A(G190), .B(new_n258), .C1(new_n274), .C2(new_n256), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n294), .A2(new_n295), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n276), .A2(new_n297), .A3(new_n293), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT73), .B1(new_n299), .B2(KEYINPUT10), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n298), .A2(new_n300), .B1(KEYINPUT10), .B2(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n275), .A2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n275), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n292), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G97), .ZN(new_n309));
  OAI211_X1 g0109(.A(G226), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n310));
  OAI211_X1 g0110(.A(G232), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT74), .B1(new_n262), .B2(G232), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n253), .B1(new_n257), .B2(G238), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT75), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n317), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT13), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT75), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(new_n322), .A3(new_n316), .A4(new_n317), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(new_n321), .A3(G179), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT79), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(KEYINPUT75), .B2(new_n318), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT79), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G179), .A4(new_n323), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(new_n318), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT14), .A3(G169), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n325), .A2(new_n329), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n290), .A2(G68), .ZN(new_n338));
  INV_X1    g0138(.A(G13), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G1), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G20), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(KEYINPUT76), .A3(G50), .ZN(new_n344));
  OAI221_X1 g0144(.A(new_n344), .B1(new_n215), .B2(G68), .C1(new_n264), .C2(new_n279), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT76), .B1(new_n277), .B2(G50), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n286), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT77), .B(KEYINPUT11), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n286), .B(new_n348), .C1(new_n345), .C2(new_n346), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n338), .B(new_n343), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT78), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n334), .B2(G200), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n319), .A2(new_n321), .A3(G190), .A4(new_n323), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n353), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n330), .B2(new_n326), .ZN(new_n360));
  AND4_X1   g0160(.A1(new_n355), .A2(new_n359), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G20), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(G33), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n215), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n363), .B1(new_n280), .B2(new_n365), .C1(new_n279), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n286), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n290), .A2(G77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n288), .A2(new_n264), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n253), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n256), .A2(new_n251), .ZN(new_n373));
  INV_X1    g0173(.A(G244), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n270), .A2(G232), .B1(G107), .B2(new_n269), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n262), .A2(G238), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n378), .B2(new_n308), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n371), .B1(new_n379), .B2(G169), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n371), .B(KEYINPUT72), .C1(new_n379), .C2(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n303), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n371), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n379), .A2(G200), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n280), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n288), .ZN(new_n393));
  INV_X1    g0193(.A(new_n290), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n392), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n260), .A2(new_n215), .A3(new_n261), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n261), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n341), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G20), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT80), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n277), .A2(new_n403), .A3(G159), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n277), .B2(G159), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT16), .B1(new_n400), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n269), .B2(new_n215), .ZN(new_n409));
  NOR4_X1   g0209(.A1(new_n267), .A2(new_n268), .A3(new_n397), .A4(G20), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  INV_X1    g0212(.A(new_n406), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n404), .B1(new_n401), .B2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n395), .B1(new_n416), .B2(new_n286), .ZN(new_n417));
  OAI211_X1 g0217(.A(G223), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n418));
  OAI211_X1 g0218(.A(G226), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n308), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT81), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n372), .B1(new_n373), .B2(new_n233), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(KEYINPUT81), .A3(new_n308), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n253), .B1(new_n257), .B2(G232), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n422), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT18), .B1(new_n417), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n421), .A2(KEYINPUT81), .A3(new_n308), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT81), .B1(new_n421), .B2(new_n308), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n426), .B1(new_n431), .B2(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(new_n286), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n408), .B2(new_n415), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n439), .C1(new_n441), .C2(new_n395), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n425), .A2(G190), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n424), .A2(new_n444), .A3(new_n427), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n430), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n412), .B1(new_n411), .B2(new_n414), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n407), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n286), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n395), .ZN(new_n452));
  AND4_X1   g0252(.A1(KEYINPUT17), .A2(new_n448), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT17), .B1(new_n417), .B2(new_n448), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n391), .A2(new_n443), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n307), .A2(new_n354), .A3(new_n362), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(G244), .C1(new_n268), .C2(new_n267), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n374), .B1(new_n260), .B2(new_n261), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(KEYINPUT4), .ZN(new_n464));
  OAI21_X1  g0264(.A(G250), .B1(new_n267), .B2(new_n268), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n259), .B1(new_n465), .B2(KEYINPUT4), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n308), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G257), .A3(new_n256), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G274), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n467), .A2(new_n387), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G250), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n260), .B2(new_n261), .ZN(new_n480));
  OAI21_X1  g0280(.A(G1698), .B1(new_n480), .B2(new_n459), .ZN(new_n481));
  INV_X1    g0281(.A(new_n462), .ZN(new_n482));
  OAI21_X1  g0282(.A(G244), .B1(new_n267), .B2(new_n268), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n459), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n484), .A3(new_n461), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n476), .B1(new_n485), .B2(new_n308), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n478), .B1(G200), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n365), .A2(new_n264), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n398), .A2(new_n399), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G107), .ZN(new_n490));
  AND2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT83), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n207), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT6), .A2(G97), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT82), .B1(new_n499), .B2(G107), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(new_n206), .A3(KEYINPUT6), .A4(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n490), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n287), .B1(G1), .B2(new_n364), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n286), .A2(new_n508), .A3(new_n205), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n287), .A2(G97), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n340), .A2(G20), .B1(new_n250), .B2(G33), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n285), .A2(new_n214), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(G97), .A4(new_n284), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(KEYINPUT84), .C1(G97), .C2(new_n287), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n506), .A2(new_n286), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n487), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n487), .B2(new_n516), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n215), .B1(new_n309), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G87), .A2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n206), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n522), .A2(new_n524), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n265), .A2(new_n215), .A3(G68), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n286), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n286), .A2(new_n508), .ZN(new_n530));
  INV_X1    g0330(.A(new_n366), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n532), .C1(new_n287), .C2(new_n531), .ZN(new_n533));
  OAI211_X1 g0333(.A(G238), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n308), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n469), .A2(new_n539), .A3(new_n479), .ZN(new_n540));
  AOI21_X1  g0340(.A(G274), .B1(new_n539), .B2(G250), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n250), .A2(G45), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n256), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n538), .A2(G179), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n431), .B1(new_n538), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n533), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n526), .A2(new_n527), .B1(new_n284), .B2(new_n513), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n531), .A2(new_n287), .ZN(new_n549));
  INV_X1    g0349(.A(G87), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n286), .A2(new_n508), .A3(new_n550), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n538), .A2(new_n387), .A3(new_n544), .ZN(new_n553));
  AOI21_X1  g0353(.A(G200), .B1(new_n538), .B2(new_n544), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT86), .B1(new_n486), .B2(new_n303), .ZN(new_n557));
  AND4_X1   g0357(.A1(KEYINPUT86), .A2(new_n467), .A3(new_n303), .A4(new_n477), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n511), .A2(new_n515), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n215), .B1(new_n498), .B2(new_n503), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n206), .B1(new_n398), .B2(new_n399), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n561), .A2(new_n562), .A3(new_n488), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n563), .B2(new_n440), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n467), .A2(new_n477), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n431), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n556), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n520), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n206), .A2(G20), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(KEYINPUT23), .B1(G20), .B2(new_n536), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT90), .B1(new_n570), .B2(KEYINPUT23), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(KEYINPUT89), .A2(G87), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n215), .B(new_n574), .C1(new_n267), .C2(new_n268), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n265), .A2(KEYINPUT22), .A3(new_n215), .A4(new_n574), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(KEYINPUT90), .A3(KEYINPUT23), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n573), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n579), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n583), .A2(new_n571), .A3(new_n572), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT24), .A3(new_n577), .A4(new_n578), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n286), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n340), .A2(G20), .A3(new_n206), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(G107), .B2(new_n530), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n465), .C2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n308), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n474), .A2(new_n469), .B1(new_n254), .B2(new_n255), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G264), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n475), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n593), .A2(new_n308), .B1(G264), .B2(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G179), .A3(new_n475), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT91), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n586), .A2(new_n589), .B1(new_n598), .B2(new_n600), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT91), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n597), .A2(G190), .ZN(new_n607));
  AOI21_X1  g0407(.A(G200), .B1(new_n599), .B2(new_n475), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n586), .B(new_n589), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n603), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(G116), .B1(new_n286), .B2(new_n508), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n287), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(G20), .B1(G33), .B2(G283), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n364), .A2(G97), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n612), .A2(G20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n286), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n286), .A2(new_n622), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n462), .B(new_n215), .C1(G33), .C2(new_n205), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n618), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT20), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n614), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  INV_X1    g0432(.A(new_n471), .ZN(new_n633));
  NAND2_X1  g0433(.A1(KEYINPUT5), .A2(G41), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n542), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n595), .A2(G270), .B1(G274), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n637));
  OAI211_X1 g0437(.A(G257), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n260), .A2(G303), .A3(new_n261), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n308), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n632), .B(new_n431), .C1(new_n636), .C2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n636), .A2(G179), .A3(new_n641), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n631), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n624), .B1(new_n621), .B2(new_n623), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n626), .A2(KEYINPUT20), .A3(new_n629), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n645), .A2(new_n646), .B1(new_n613), .B2(new_n611), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n636), .A2(new_n641), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G169), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n632), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n648), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G200), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n648), .A2(G190), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n610), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n458), .A2(new_n569), .A3(new_n657), .ZN(G372));
  AOI211_X1 g0458(.A(G190), .B(new_n476), .C1(new_n485), .C2(new_n308), .ZN(new_n659));
  AOI21_X1  g0459(.A(G200), .B1(new_n467), .B2(new_n477), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT85), .B1(new_n661), .B2(new_n564), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n487), .A2(new_n516), .A3(new_n517), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n547), .A2(new_n555), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT86), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n565), .B2(G179), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n486), .A2(KEYINPUT86), .A3(new_n303), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n506), .A2(new_n286), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n560), .B1(new_n431), .B2(new_n565), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n665), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n664), .A2(new_n672), .A3(new_n609), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n644), .A2(new_n650), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT92), .B1(new_n674), .B2(new_n604), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n602), .A2(new_n676), .A3(new_n650), .A4(new_n644), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n559), .A2(new_n567), .ZN(new_n680));
  XOR2_X1   g0480(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n556), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n669), .A2(new_n671), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n665), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n682), .B(new_n547), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n458), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n356), .A2(new_n357), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n383), .A3(new_n382), .A4(new_n384), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n354), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT17), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n448), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n443), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n298), .A2(new_n300), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n306), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n701), .ZN(G369));
  INV_X1    g0502(.A(new_n340), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .A3(G20), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT27), .B1(new_n703), .B2(G20), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n647), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n656), .B2(KEYINPUT94), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n655), .A2(new_n650), .A3(new_n644), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT94), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n712), .A2(new_n715), .B1(new_n651), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n590), .A2(new_n708), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n603), .A2(new_n606), .A3(new_n609), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n604), .A2(new_n708), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n716), .A2(G330), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n674), .A2(new_n709), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n718), .A2(new_n722), .B1(new_n602), .B2(new_n708), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(G399));
  NAND3_X1  g0525(.A1(new_n523), .A2(new_n206), .A3(new_n612), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT95), .Z(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n250), .ZN(new_n728));
  INV_X1    g0528(.A(new_n211), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  MUX2_X1   g0530(.A(new_n728), .B(new_n218), .S(new_n730), .Z(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n684), .A2(new_n685), .ZN(new_n733));
  INV_X1    g0533(.A(new_n681), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n683), .B2(new_n665), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n547), .B(KEYINPUT97), .Z(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT98), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n664), .A2(new_n672), .A3(new_n609), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n651), .A2(new_n603), .A3(new_n606), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n590), .A2(new_n601), .A3(new_n605), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n605), .B1(new_n590), .B2(new_n601), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n743), .A2(new_n744), .A3(new_n674), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n673), .A2(new_n745), .A3(KEYINPUT98), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n738), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT99), .B1(new_n747), .B2(new_n709), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n569), .A2(new_n739), .A3(new_n609), .A4(new_n741), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT98), .B1(new_n673), .B2(new_n745), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n737), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT99), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n751), .A2(new_n752), .A3(new_n708), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT29), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n687), .A2(new_n709), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n486), .A2(new_n544), .A3(new_n538), .A4(new_n599), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  INV_X1    g0559(.A(new_n643), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(new_n762));
  AOI21_X1  g0562(.A(G179), .B1(new_n538), .B2(new_n544), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n565), .A2(new_n597), .A3(new_n648), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(new_n766), .A3(new_n708), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n657), .A2(new_n569), .A3(new_n709), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(new_n765), .B2(new_n708), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT96), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(KEYINPUT96), .A3(G330), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n757), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n732), .B1(new_n778), .B2(G1), .ZN(G364));
  NOR2_X1   g0579(.A1(new_n339), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n250), .B1(new_n780), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n730), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n211), .A2(new_n265), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G355), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G116), .B2(new_n211), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT101), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n729), .A2(new_n265), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n248), .A2(new_n468), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n218), .A2(G45), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n214), .B1(G20), .B2(new_n431), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n215), .A2(new_n387), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n803), .A2(new_n446), .A3(G179), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n215), .A2(G190), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(G179), .A3(new_n446), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n805), .A2(new_n550), .B1(new_n809), .B2(new_n206), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n303), .A2(new_n446), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n269), .B(new_n810), .C1(G50), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G179), .A2(G200), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n215), .B1(new_n815), .B2(G190), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G97), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n806), .A2(new_n815), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n803), .A2(new_n303), .A3(G200), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G58), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n811), .A2(new_n806), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n341), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n807), .A2(new_n303), .A3(G200), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(G77), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n814), .A2(new_n821), .A3(new_n825), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G322), .ZN(new_n834));
  INV_X1    g0634(.A(G326), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n827), .A2(new_n834), .B1(new_n812), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n265), .B(new_n836), .C1(G311), .C2(new_n831), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n820), .A2(G294), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n822), .B(KEYINPUT103), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G329), .ZN(new_n840));
  INV_X1    g0640(.A(new_n829), .ZN(new_n841));
  NOR2_X1   g0641(.A1(KEYINPUT33), .A2(G317), .ZN(new_n842));
  AND2_X1   g0642(.A1(KEYINPUT33), .A2(G317), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n809), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G303), .B2(new_n804), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n837), .A2(new_n838), .A3(new_n840), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n784), .B(new_n801), .C1(new_n799), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n798), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n716), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n783), .B1(new_n716), .B2(G330), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(G330), .B2(new_n716), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  NOR2_X1   g0656(.A1(new_n386), .A2(new_n709), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n385), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n385), .B2(new_n390), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT106), .ZN(new_n862));
  MUX2_X1   g0662(.A(new_n862), .B(new_n861), .S(new_n755), .Z(new_n863));
  OR2_X1    g0663(.A1(new_n863), .A2(new_n776), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n776), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n784), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n799), .A2(new_n796), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n783), .B1(G77), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(G303), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n809), .A2(new_n550), .B1(new_n870), .B2(new_n812), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n265), .B(new_n871), .C1(G283), .C2(new_n841), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n839), .A2(G311), .ZN(new_n873));
  INV_X1    g0673(.A(G294), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n206), .A2(new_n805), .B1(new_n827), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G116), .B2(new_n831), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n821), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G50), .A2(new_n804), .B1(new_n808), .B2(G68), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT104), .Z(new_n879));
  AOI22_X1  g0679(.A1(new_n831), .A2(G159), .B1(new_n813), .B2(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  INV_X1    g0681(.A(G143), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n881), .B2(new_n829), .C1(new_n882), .C2(new_n827), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT34), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n879), .B(new_n885), .C1(new_n828), .C2(new_n819), .ZN(new_n886));
  INV_X1    g0686(.A(G132), .ZN(new_n887));
  INV_X1    g0687(.A(new_n839), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n265), .B1(new_n887), .B2(new_n888), .C1(new_n883), .C2(new_n884), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n877), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n869), .B1(new_n890), .B2(new_n799), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT105), .Z(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n797), .B2(new_n861), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n866), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(new_n701), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT29), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n747), .A2(KEYINPUT99), .A3(new_n709), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n752), .B1(new_n751), .B2(new_n708), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n755), .A2(KEYINPUT29), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n895), .B1(new_n901), .B2(new_n458), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT109), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n336), .B1(new_n358), .B2(new_n361), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n353), .A2(new_n708), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n689), .B(new_n905), .C1(new_n336), .C2(new_n359), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n709), .B(new_n861), .C1(new_n679), .C2(new_n686), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n385), .A2(new_n708), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT107), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT108), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n910), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(new_n706), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n441), .B2(new_n395), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n443), .B2(new_n455), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n428), .B(new_n432), .C1(new_n441), .C2(new_n395), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n692), .A3(new_n921), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT37), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n923), .A2(new_n692), .A3(KEYINPUT37), .A4(new_n921), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n919), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n434), .A2(new_n442), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n696), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(KEYINPUT38), .A3(new_n926), .A4(new_n927), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(KEYINPUT39), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n354), .A2(new_n708), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n936), .A2(new_n937), .B1(new_n931), .B2(new_n706), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n903), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n858), .B1(new_n391), .B2(new_n857), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n907), .B2(new_n908), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n771), .A3(new_n934), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(KEYINPUT110), .A3(KEYINPUT40), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n771), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n457), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G330), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n940), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n940), .A2(new_n953), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n250), .C2(new_n780), .ZN(new_n956));
  OAI21_X1  g0756(.A(G77), .B1(new_n828), .B2(new_n341), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n957), .A2(new_n217), .B1(G50), .B2(new_n341), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(G1), .A3(new_n339), .ZN(new_n959));
  OAI211_X1 g0759(.A(G116), .B(new_n216), .C1(new_n504), .C2(KEYINPUT35), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(KEYINPUT35), .B2(new_n504), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT36), .Z(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT111), .ZN(G367));
  AND2_X1   g0764(.A1(new_n239), .A2(new_n791), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n800), .B1(new_n211), .B2(new_n366), .ZN(new_n966));
  INV_X1    g0766(.A(new_n831), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n202), .A2(new_n967), .B1(new_n809), .B2(new_n264), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n827), .A2(new_n881), .B1(new_n829), .B2(new_n823), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n820), .A2(G68), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n269), .B1(new_n813), .B2(G143), .ZN(new_n972));
  INV_X1    g0772(.A(new_n822), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n804), .A2(G58), .B1(G137), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n809), .A2(new_n205), .B1(new_n874), .B2(new_n829), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n265), .B(new_n976), .C1(G311), .C2(new_n813), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n804), .A2(G116), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n831), .A2(G283), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n826), .A2(G303), .B1(G317), .B2(new_n973), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n819), .A2(new_n206), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT47), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n799), .B1(new_n984), .B2(new_n985), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n783), .B1(new_n965), .B2(new_n966), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT114), .Z(new_n989));
  OR2_X1    g0789(.A1(new_n709), .A2(new_n552), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n556), .A2(KEYINPUT112), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n547), .B2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT112), .B1(new_n556), .B2(new_n990), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n989), .B1(new_n851), .B2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n669), .A2(new_n671), .B1(new_n564), .B2(new_n708), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n664), .A2(new_n997), .B1(new_n680), .B2(new_n708), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n998), .A2(new_n718), .A3(new_n722), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n664), .A2(new_n997), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n743), .A2(new_n744), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n683), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n709), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1000), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n994), .A2(KEYINPUT113), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1009), .B1(KEYINPUT43), .B2(new_n995), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n721), .A2(new_n998), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n723), .A2(new_n998), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT44), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n998), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n724), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n723), .B2(new_n998), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1018), .A2(new_n721), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n656), .A2(KEYINPUT94), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n1026), .B1(new_n674), .B2(new_n710), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n720), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1027), .A2(new_n952), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1023), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n1017), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1028), .B1(new_n1027), .B2(new_n952), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n722), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n1033), .A2(new_n721), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1033), .B2(new_n721), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n757), .B(new_n776), .C1(new_n1032), .C2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n730), .B(KEYINPUT41), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n782), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n996), .B1(new_n1015), .B2(new_n1042), .ZN(G387));
  OAI211_X1 g0843(.A(new_n1037), .B(new_n776), .C1(new_n899), .C2(new_n900), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n730), .ZN(new_n1046));
  OAI21_X1  g0846(.A(KEYINPUT116), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT116), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1044), .A2(new_n1048), .A3(new_n730), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n777), .A2(new_n1038), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1028), .A2(new_n798), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n786), .A2(new_n727), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(G107), .B2(new_n211), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n234), .A2(G45), .ZN(new_n1055));
  AOI211_X1 g0855(.A(G45), .B(new_n727), .C1(G68), .C2(G77), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n280), .A2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n729), .B(new_n265), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1054), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n800), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n783), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n805), .A2(new_n264), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n265), .B1(new_n809), .B2(new_n205), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G159), .C2(new_n813), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n820), .A2(new_n531), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n826), .A2(G50), .B1(G150), .B2(new_n973), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n831), .A2(G68), .B1(new_n841), .B2(new_n392), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G322), .A2(new_n813), .B1(new_n841), .B2(G311), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT115), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G317), .A2(new_n826), .B1(new_n831), .B2(G303), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n819), .A2(new_n845), .B1(new_n805), .B2(new_n874), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1074), .B2(KEYINPUT48), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n265), .B1(new_n808), .B2(G116), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n835), .C2(new_n822), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT49), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1069), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1062), .B1(new_n1082), .B2(new_n799), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1037), .A2(new_n782), .B1(new_n1052), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1051), .A2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n1032), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1046), .B1(new_n1045), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1045), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n244), .A2(new_n729), .A3(new_n265), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n800), .B1(new_n211), .B2(new_n205), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n805), .A2(new_n845), .B1(new_n967), .B2(new_n874), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n829), .A2(new_n870), .B1(new_n822), .B2(new_n834), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n265), .B1(new_n808), .B2(G107), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(new_n612), .C2(new_n819), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n826), .A2(G311), .B1(new_n813), .B2(G317), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n805), .A2(new_n341), .B1(new_n967), .B2(new_n280), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n829), .A2(new_n202), .B1(new_n822), .B2(new_n882), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n820), .A2(G77), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n269), .B1(new_n808), .B2(G87), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n826), .A2(G159), .B1(new_n813), .B2(G150), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1095), .A2(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n799), .B1(new_n1107), .B2(KEYINPUT118), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n783), .B1(new_n1089), .B2(new_n1090), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n798), .B2(new_n998), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1086), .B2(new_n782), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1088), .A2(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n936), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n796), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n783), .B1(new_n392), .B2(new_n868), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n809), .A2(new_n341), .B1(new_n206), .B2(new_n829), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n265), .B(new_n1117), .C1(G87), .C2(new_n804), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n839), .A2(G294), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n827), .A2(new_n612), .B1(new_n812), .B2(new_n845), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G97), .B2(new_n831), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1102), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n819), .A2(new_n823), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n827), .A2(new_n887), .B1(new_n812), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G137), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n809), .A2(new_n202), .B1(new_n1126), .B2(new_n829), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n804), .A2(G150), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n269), .B1(new_n831), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n839), .A2(G125), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1128), .A2(new_n1131), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1122), .B1(new_n1123), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1116), .B1(new_n1137), .B2(new_n799), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1115), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1114), .B1(new_n918), .B2(new_n937), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n774), .A2(new_n775), .A3(new_n942), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n861), .B1(new_n748), .B2(new_n753), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n912), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n910), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n937), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n934), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1140), .B(new_n1141), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n915), .A2(new_n917), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1148), .B2(new_n910), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n941), .B1(new_n897), .B2(new_n898), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n909), .B1(new_n1150), .B2(new_n912), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1146), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1149), .A2(new_n1114), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n772), .A2(new_n910), .A3(new_n941), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1147), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1139), .B1(new_n1156), .B2(new_n781), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n754), .A2(new_n756), .A3(new_n458), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n950), .A2(G330), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n701), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT119), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT119), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .A4(new_n701), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n774), .A2(new_n775), .A3(new_n861), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1154), .B1(new_n1165), .B2(new_n910), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n910), .B1(new_n772), .B2(new_n862), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1141), .A2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1166), .A2(new_n1148), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1162), .A2(new_n1164), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1147), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1155), .B1(new_n1174), .B2(new_n1140), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n730), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1171), .A2(new_n1156), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1158), .B1(new_n1177), .B2(new_n1178), .ZN(G378));
  AOI21_X1  g0979(.A(new_n784), .B1(new_n202), .B2(new_n867), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n804), .A2(new_n1133), .B1(G132), .B2(new_n841), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1124), .B2(new_n827), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n831), .A2(G137), .B1(new_n813), .B2(G125), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n881), .C2(new_n819), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  INV_X1    g0987(.A(G41), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n364), .B(new_n1188), .C1(new_n809), .C2(new_n823), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G124), .B2(new_n973), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n826), .A2(G107), .B1(new_n813), .B2(G116), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n205), .B2(new_n829), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n366), .A2(new_n967), .B1(new_n809), .B2(new_n828), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n269), .A2(new_n1188), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1063), .A4(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n971), .C1(new_n845), .C2(new_n888), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1195), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1201));
  AND4_X1   g1001(.A1(new_n1191), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT121), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n799), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n292), .A2(new_n920), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n307), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1206), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n301), .B2(new_n306), .ZN(new_n1209));
  XOR2_X1   g1009(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1207), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1206), .B1(new_n700), .B2(new_n305), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n301), .A2(new_n306), .A3(new_n1208), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1210), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1180), .B1(new_n1203), .B2(new_n1205), .C1(new_n1216), .C2(new_n797), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n943), .A2(KEYINPUT110), .A3(KEYINPUT40), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT40), .B1(new_n943), .B2(KEYINPUT110), .ZN(new_n1220));
  OAI21_X1  g1020(.A(G330), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G330), .B(new_n1216), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n935), .A3(new_n938), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1216), .B1(new_n948), .B2(G330), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1223), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n939), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1218), .B1(new_n1228), .B2(new_n782), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT122), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1230), .B(new_n939), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1224), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1230), .B1(new_n1233), .B2(new_n939), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1176), .B2(new_n1170), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n730), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1170), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1164), .B(new_n1162), .C1(new_n1156), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1228), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1229), .B1(new_n1238), .B2(new_n1241), .ZN(G375));
  AOI21_X1  g1042(.A(new_n1163), .B1(new_n902), .B2(new_n1160), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1164), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1239), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n1041), .A3(new_n1171), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n910), .A2(new_n796), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n783), .B1(G68), .B2(new_n868), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT123), .Z(new_n1249));
  OAI22_X1  g1049(.A1(new_n827), .A2(new_n845), .B1(new_n967), .B2(new_n206), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n265), .B(new_n1250), .C1(G77), .C2(new_n808), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n839), .A2(G303), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n805), .A2(new_n205), .B1(new_n829), .B2(new_n612), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G294), .B2(new_n813), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(new_n1066), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n265), .B1(new_n809), .B2(new_n828), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n1124), .C2(new_n888), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1126), .A2(new_n827), .B1(new_n805), .B2(new_n823), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G150), .B2(new_n831), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n813), .A2(G132), .B1(new_n841), .B2(new_n1133), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n202), .C2(new_n819), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1255), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1249), .B1(new_n799), .B2(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1170), .A2(new_n782), .B1(new_n1247), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(new_n1178), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1046), .B1(new_n1171), .B2(new_n1156), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1157), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1270), .B(new_n1229), .C1(new_n1238), .C2(new_n1241), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1051), .A2(new_n855), .A3(new_n1084), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(G390), .A2(new_n1273), .A3(G387), .A4(G384), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1272), .A2(new_n1266), .A3(new_n1246), .A4(new_n1274), .ZN(G407));
  OAI211_X1 g1075(.A(G407), .B(G213), .C1(G343), .C2(new_n1271), .ZN(G409));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G387), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1273), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n855), .B1(new_n1051), .B2(new_n1084), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(G387), .A3(new_n1273), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1281), .A2(G390), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G390), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1229), .C1(new_n1238), .C2(new_n1241), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1228), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1237), .A2(new_n1040), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n782), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1217), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1270), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n707), .A2(G213), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1171), .A2(new_n730), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1245), .A2(KEYINPUT60), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1236), .A2(new_n1298), .A3(new_n1239), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(G384), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1266), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1296), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1298), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1305));
  AOI211_X1 g1105(.A(KEYINPUT60), .B(new_n1170), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G384), .B1(new_n1307), .B2(new_n1266), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1303), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .A4(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT61), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1287), .A2(new_n1292), .B1(G213), .B2(new_n707), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n707), .A2(G213), .A3(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1301), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1307), .A2(G384), .A3(new_n1266), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1313), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1310), .B(new_n1311), .C1(new_n1312), .C2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1294), .B1(new_n1312), .B2(new_n1309), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1286), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1311), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1295), .A4(new_n1309), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT126), .B(new_n1311), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT63), .B1(new_n1319), .B2(new_n1312), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1312), .A2(new_n1309), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1322), .A2(new_n1332), .ZN(G405));
  INV_X1    g1133(.A(KEYINPUT57), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1237), .B2(new_n1288), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1227), .A2(KEYINPUT122), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(new_n1224), .A3(new_n1231), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1337), .A2(new_n1240), .A3(KEYINPUT57), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1335), .A2(new_n730), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1270), .B1(new_n1339), .B2(new_n1229), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1309), .B1(new_n1272), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1286), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G375), .A2(G378), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1271), .A3(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(new_n1342), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1342), .B1(new_n1341), .B2(new_n1345), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1346), .B1(new_n1347), .B2(KEYINPUT127), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT127), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1349), .B(new_n1342), .C1(new_n1341), .C2(new_n1345), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(G402));
endmodule


