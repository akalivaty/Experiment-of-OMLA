

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U548 ( .A1(n676), .A2(n769), .ZN(n714) );
  XNOR2_X1 U549 ( .A(n576), .B(KEYINPUT71), .ZN(n578) );
  NAND2_X2 U550 ( .A1(n578), .A2(n577), .ZN(n1003) );
  NOR2_X2 U551 ( .A1(G164), .A2(G1384), .ZN(n770) );
  NOR2_X1 U552 ( .A1(n694), .A2(n693), .ZN(n695) );
  BUF_X1 U553 ( .A(n549), .Z(n533) );
  AND2_X1 U554 ( .A1(n698), .A2(n512), .ZN(n699) );
  XNOR2_X1 U555 ( .A(KEYINPUT28), .B(n697), .ZN(n512) );
  NOR2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n513) );
  NOR2_X1 U557 ( .A1(G651), .A2(n624), .ZN(n638) );
  XOR2_X2 U558 ( .A(n513), .B(KEYINPUT17), .Z(n978) );
  NAND2_X1 U559 ( .A1(G138), .A2(n978), .ZN(n515) );
  XOR2_X1 U560 ( .A(KEYINPUT64), .B(G2104), .Z(n516) );
  AND2_X1 U561 ( .A1(n516), .A2(G2105), .ZN(n975) );
  NAND2_X1 U562 ( .A1(G126), .A2(n975), .ZN(n514) );
  NAND2_X1 U563 ( .A1(n515), .A2(n514), .ZN(n520) );
  AND2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n976) );
  NAND2_X1 U565 ( .A1(G114), .A2(n976), .ZN(n518) );
  NOR2_X1 U566 ( .A1(n516), .A2(G2105), .ZN(n549) );
  NAND2_X1 U567 ( .A1(G102), .A2(n549), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U569 ( .A1(n520), .A2(n519), .ZN(G164) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n630) );
  NAND2_X1 U571 ( .A1(G85), .A2(n630), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n624) );
  INV_X1 U573 ( .A(G651), .ZN(n523) );
  NOR2_X1 U574 ( .A1(n624), .A2(n523), .ZN(n634) );
  NAND2_X1 U575 ( .A1(G72), .A2(n634), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n524), .Z(n631) );
  NAND2_X1 U579 ( .A1(G60), .A2(n631), .ZN(n526) );
  NAND2_X1 U580 ( .A1(G47), .A2(n638), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U582 ( .A1(n528), .A2(n527), .ZN(G290) );
  XNOR2_X1 U583 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U584 ( .A1(n975), .A2(G123), .ZN(n530) );
  XNOR2_X1 U585 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n530), .B(n529), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G135), .A2(n978), .ZN(n532) );
  NAND2_X1 U588 ( .A1(G111), .A2(n976), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G99), .A2(n533), .ZN(n534) );
  XNOR2_X1 U591 ( .A(KEYINPUT75), .B(n534), .ZN(n535) );
  NOR2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n987) );
  XNOR2_X1 U594 ( .A(G2096), .B(n987), .ZN(n539) );
  OR2_X1 U595 ( .A1(G2100), .A2(n539), .ZN(G156) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  INV_X1 U598 ( .A(G120), .ZN(G236) );
  INV_X1 U599 ( .A(G69), .ZN(G235) );
  INV_X1 U600 ( .A(G108), .ZN(G238) );
  NAND2_X1 U601 ( .A1(n638), .A2(G52), .ZN(n540) );
  XNOR2_X1 U602 ( .A(KEYINPUT65), .B(n540), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G90), .A2(n630), .ZN(n542) );
  NAND2_X1 U604 ( .A1(G77), .A2(n634), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n543), .B(KEYINPUT9), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT66), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n631), .A2(G64), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(G171) );
  INV_X1 U611 ( .A(G171), .ZN(G301) );
  NAND2_X1 U612 ( .A1(n976), .A2(G113), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G101), .A2(n549), .ZN(n550) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n550), .Z(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n673) );
  NAND2_X1 U616 ( .A1(G125), .A2(n975), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G137), .A2(n978), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n671) );
  NOR2_X1 U619 ( .A1(n673), .A2(n671), .ZN(G160) );
  NAND2_X1 U620 ( .A1(n630), .A2(G89), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G76), .A2(n634), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G63), .A2(n631), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G51), .A2(n638), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G94), .A2(G452), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n566) );
  XOR2_X1 U635 ( .A(n566), .B(KEYINPUT10), .Z(n1016) );
  NAND2_X1 U636 ( .A1(n1016), .A2(G567), .ZN(n567) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U638 ( .A1(n630), .A2(G81), .ZN(n568) );
  XNOR2_X1 U639 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G68), .A2(n634), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U642 ( .A(n571), .B(KEYINPUT13), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G56), .A2(n631), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT70), .ZN(n573) );
  XNOR2_X1 U645 ( .A(KEYINPUT14), .B(n573), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U647 ( .A1(G43), .A2(n638), .ZN(n577) );
  INV_X1 U648 ( .A(G860), .ZN(n600) );
  OR2_X1 U649 ( .A1(n1003), .A2(n600), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U651 ( .A1(G92), .A2(n630), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G79), .A2(n634), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G66), .A2(n631), .ZN(n582) );
  NAND2_X1 U655 ( .A1(G54), .A2(n638), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n585), .Z(n1004) );
  OR2_X1 U659 ( .A1(n1004), .A2(G868), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G91), .A2(n630), .ZN(n588) );
  XOR2_X1 U662 ( .A(KEYINPUT68), .B(n588), .Z(n593) );
  NAND2_X1 U663 ( .A1(G65), .A2(n631), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G53), .A2(n638), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U666 ( .A(KEYINPUT69), .B(n591), .Z(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n634), .A2(G78), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G299) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT72), .ZN(n598) );
  INV_X1 U672 ( .A(G868), .ZN(n650) );
  NOR2_X1 U673 ( .A1(n650), .A2(G286), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U675 ( .A(KEYINPUT73), .B(n599), .Z(G297) );
  NAND2_X1 U676 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n601), .A2(n1004), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n1003), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G868), .A2(n1004), .ZN(n603) );
  NOR2_X1 U681 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G93), .A2(n630), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G80), .A2(n634), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G67), .A2(n631), .ZN(n608) );
  XNOR2_X1 U687 ( .A(KEYINPUT77), .B(n608), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n638), .A2(G55), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n649) );
  XNOR2_X1 U691 ( .A(n1003), .B(KEYINPUT76), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n1004), .A2(G559), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n614), .B(n613), .ZN(n646) );
  NOR2_X1 U694 ( .A1(n646), .A2(G860), .ZN(n615) );
  XOR2_X1 U695 ( .A(n649), .B(n615), .Z(G145) );
  NAND2_X1 U696 ( .A1(G75), .A2(n634), .ZN(n617) );
  NAND2_X1 U697 ( .A1(G62), .A2(n631), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G88), .A2(n630), .ZN(n618) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n618), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n638), .A2(G50), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(G303) );
  NAND2_X1 U704 ( .A1(G49), .A2(n638), .ZN(n623) );
  XNOR2_X1 U705 ( .A(n623), .B(KEYINPUT78), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G87), .A2(n624), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n631), .A2(n627), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G86), .A2(n630), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G61), .A2(n631), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n634), .A2(G73), .ZN(n635) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n638), .A2(G48), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(G305) );
  XOR2_X1 U719 ( .A(G303), .B(KEYINPUT19), .Z(n645) );
  XNOR2_X1 U720 ( .A(G290), .B(G288), .ZN(n643) );
  XNOR2_X1 U721 ( .A(G299), .B(G305), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n641), .B(n649), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n645), .B(n644), .ZN(n1007) );
  XNOR2_X1 U725 ( .A(n646), .B(n1007), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n647), .A2(G868), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT80), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U730 ( .A1(G2084), .A2(G2078), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(KEYINPUT20), .ZN(n654) );
  XNOR2_X1 U732 ( .A(KEYINPUT81), .B(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n655), .A2(G2090), .ZN(n656) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(n656), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(G2072), .ZN(G158) );
  NOR2_X1 U736 ( .A1(G235), .A2(G236), .ZN(n658) );
  XOR2_X1 U737 ( .A(KEYINPUT82), .B(n658), .Z(n659) );
  NOR2_X1 U738 ( .A1(G238), .A2(n659), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G57), .A2(n660), .ZN(n951) );
  NAND2_X1 U740 ( .A1(G567), .A2(n951), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n661), .B(KEYINPUT83), .ZN(n666) );
  NOR2_X1 U742 ( .A1(G220), .A2(G219), .ZN(n662) );
  XNOR2_X1 U743 ( .A(KEYINPUT22), .B(n662), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n663), .A2(G96), .ZN(n664) );
  OR2_X1 U745 ( .A1(G218), .A2(n664), .ZN(n952) );
  AND2_X1 U746 ( .A1(G2106), .A2(n952), .ZN(n665) );
  NOR2_X1 U747 ( .A1(n666), .A2(n665), .ZN(G319) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n668) );
  INV_X1 U749 ( .A(G319), .ZN(n667) );
  NOR2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U751 ( .A(n669), .B(KEYINPUT84), .ZN(n832) );
  NAND2_X1 U752 ( .A1(G36), .A2(n832), .ZN(G176) );
  INV_X1 U753 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U754 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n700) );
  INV_X1 U755 ( .A(n770), .ZN(n676) );
  INV_X1 U756 ( .A(G40), .ZN(n670) );
  OR2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n769) );
  NOR2_X1 U759 ( .A1(n676), .A2(n769), .ZN(n674) );
  NAND2_X1 U760 ( .A1(G1996), .A2(n674), .ZN(n675) );
  XNOR2_X1 U761 ( .A(n675), .B(KEYINPUT26), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G1341), .A2(n714), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U764 ( .A(KEYINPUT93), .B(n679), .Z(n680) );
  NOR2_X2 U765 ( .A1(n680), .A2(n1003), .ZN(n681) );
  OR2_X1 U766 ( .A1(n1004), .A2(n681), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n681), .A2(n1004), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G1348), .A2(n714), .ZN(n683) );
  XOR2_X1 U769 ( .A(n714), .B(KEYINPUT92), .Z(n701) );
  NAND2_X1 U770 ( .A1(G2067), .A2(n701), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U774 ( .A(KEYINPUT94), .B(n688), .Z(n694) );
  NAND2_X1 U775 ( .A1(G2072), .A2(n701), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT27), .B(n689), .Z(n692) );
  INV_X1 U777 ( .A(n701), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n690), .A2(G1956), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U780 ( .A1(G299), .A2(n696), .ZN(n693) );
  XNOR2_X1 U781 ( .A(n695), .B(KEYINPUT95), .ZN(n698) );
  NAND2_X1 U782 ( .A1(G299), .A2(n696), .ZN(n697) );
  XNOR2_X1 U783 ( .A(n700), .B(n699), .ZN(n727) );
  XNOR2_X1 U784 ( .A(G2078), .B(KEYINPUT25), .ZN(n850) );
  NAND2_X1 U785 ( .A1(n701), .A2(n850), .ZN(n703) );
  INV_X1 U786 ( .A(G1961), .ZN(n953) );
  NAND2_X1 U787 ( .A1(n953), .A2(n714), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n708) );
  NAND2_X1 U789 ( .A1(G171), .A2(n708), .ZN(n726) );
  AND2_X1 U790 ( .A1(n726), .A2(G286), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n727), .A2(n704), .ZN(n721) );
  INV_X1 U792 ( .A(G286), .ZN(n713) );
  NAND2_X1 U793 ( .A1(G8), .A2(n714), .ZN(n765) );
  NOR2_X1 U794 ( .A1(G1966), .A2(n765), .ZN(n731) );
  NOR2_X1 U795 ( .A1(G2084), .A2(n714), .ZN(n725) );
  NOR2_X1 U796 ( .A1(n731), .A2(n725), .ZN(n705) );
  NAND2_X1 U797 ( .A1(G8), .A2(n705), .ZN(n706) );
  XNOR2_X1 U798 ( .A(KEYINPUT30), .B(n706), .ZN(n707) );
  NOR2_X1 U799 ( .A1(G168), .A2(n707), .ZN(n710) );
  NOR2_X1 U800 ( .A1(G171), .A2(n708), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U802 ( .A(KEYINPUT97), .B(n711), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n712), .B(KEYINPUT31), .ZN(n729) );
  OR2_X1 U804 ( .A1(n713), .A2(n729), .ZN(n719) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n765), .ZN(n716) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n714), .ZN(n715) );
  NOR2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n717), .A2(G303), .ZN(n718) );
  AND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n722), .B(KEYINPUT98), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n723), .A2(G8), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n724), .B(KEYINPUT32), .ZN(n735) );
  NAND2_X1 U814 ( .A1(G8), .A2(n725), .ZN(n733) );
  NAND2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n728) );
  AND2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U819 ( .A1(n735), .A2(n734), .ZN(n762) );
  INV_X1 U820 ( .A(n762), .ZN(n738) );
  NOR2_X1 U821 ( .A1(G1976), .A2(G288), .ZN(n740) );
  NOR2_X1 U822 ( .A1(G1971), .A2(G303), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n740), .A2(n736), .ZN(n869) );
  XNOR2_X1 U824 ( .A(KEYINPUT99), .B(n869), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U826 ( .A1(n739), .A2(n765), .ZN(n747) );
  NAND2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n865) );
  INV_X1 U828 ( .A(KEYINPUT33), .ZN(n749) );
  INV_X1 U829 ( .A(n765), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n749), .A2(n742), .ZN(n743) );
  XOR2_X1 U832 ( .A(n743), .B(KEYINPUT100), .Z(n748) );
  AND2_X1 U833 ( .A1(n865), .A2(n748), .ZN(n745) );
  XNOR2_X1 U834 ( .A(G1981), .B(G305), .ZN(n860) );
  INV_X1 U835 ( .A(n860), .ZN(n744) );
  AND2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n758) );
  INV_X1 U838 ( .A(n748), .ZN(n750) );
  OR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n860), .A2(n751), .ZN(n756) );
  NOR2_X1 U841 ( .A1(G1981), .A2(G305), .ZN(n752) );
  XNOR2_X1 U842 ( .A(n752), .B(KEYINPUT91), .ZN(n753) );
  XNOR2_X1 U843 ( .A(n753), .B(KEYINPUT24), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n754), .A2(n765), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  AND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n767) );
  NAND2_X1 U847 ( .A1(G8), .A2(G166), .ZN(n759) );
  NOR2_X1 U848 ( .A1(G2090), .A2(n759), .ZN(n760) );
  XNOR2_X1 U849 ( .A(n760), .B(KEYINPUT101), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(KEYINPUT102), .B(n763), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n803) );
  XOR2_X1 U854 ( .A(G1986), .B(KEYINPUT85), .Z(n768) );
  XNOR2_X1 U855 ( .A(G290), .B(n768), .ZN(n871) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n814) );
  NAND2_X1 U857 ( .A1(n871), .A2(n814), .ZN(n801) );
  NAND2_X1 U858 ( .A1(G141), .A2(n978), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G117), .A2(n976), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n533), .A2(G105), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT38), .B(n773), .Z(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n975), .A2(G129), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n993) );
  NAND2_X1 U866 ( .A1(G1996), .A2(n993), .ZN(n785) );
  NAND2_X1 U867 ( .A1(G119), .A2(n975), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G107), .A2(n976), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G131), .A2(n978), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G95), .A2(n533), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n990) );
  NAND2_X1 U874 ( .A1(G1991), .A2(n990), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n932) );
  NAND2_X1 U876 ( .A1(n932), .A2(n814), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT89), .ZN(n807) );
  XOR2_X1 U878 ( .A(KEYINPUT90), .B(n807), .Z(n799) );
  NAND2_X1 U879 ( .A1(G140), .A2(n978), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G104), .A2(n533), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n790) );
  XOR2_X1 U882 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n789) );
  XNOR2_X1 U883 ( .A(n790), .B(n789), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G128), .A2(n975), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G116), .A2(n976), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT36), .ZN(n797) );
  XNOR2_X1 U890 ( .A(n797), .B(KEYINPUT88), .ZN(n1001) );
  XNOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .ZN(n798) );
  XNOR2_X1 U892 ( .A(n798), .B(KEYINPUT86), .ZN(n812) );
  NOR2_X1 U893 ( .A1(n1001), .A2(n812), .ZN(n929) );
  NAND2_X1 U894 ( .A1(n814), .A2(n929), .ZN(n810) );
  AND2_X1 U895 ( .A1(n799), .A2(n810), .ZN(n800) );
  AND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n993), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT103), .B(n804), .Z(n937) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n990), .ZN(n926) );
  NOR2_X1 U902 ( .A1(n805), .A2(n926), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n937), .A2(n808), .ZN(n809) );
  XNOR2_X1 U905 ( .A(KEYINPUT39), .B(n809), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n1001), .A2(n812), .ZN(n933) );
  NAND2_X1 U908 ( .A1(n813), .A2(n933), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U912 ( .A(G1348), .B(G2454), .ZN(n819) );
  XNOR2_X1 U913 ( .A(n819), .B(G2430), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(G1341), .ZN(n826) );
  XOR2_X1 U915 ( .A(G2443), .B(G2427), .Z(n822) );
  XNOR2_X1 U916 ( .A(G2438), .B(G2446), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n822), .B(n821), .ZN(n824) );
  XOR2_X1 U918 ( .A(G2451), .B(G2435), .Z(n823) );
  XNOR2_X1 U919 ( .A(n824), .B(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n826), .B(n825), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(G14), .ZN(n1010) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(n1010), .Z(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n1016), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n829) );
  INV_X1 U925 ( .A(G661), .ZN(n828) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n830), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U930 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NAND2_X1 U932 ( .A1(G136), .A2(n978), .ZN(n834) );
  NAND2_X1 U933 ( .A1(G112), .A2(n976), .ZN(n833) );
  NAND2_X1 U934 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n975), .A2(G124), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n835), .B(KEYINPUT44), .ZN(n837) );
  NAND2_X1 U937 ( .A1(G100), .A2(n533), .ZN(n836) );
  NAND2_X1 U938 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U939 ( .A1(n839), .A2(n838), .ZN(G162) );
  XOR2_X1 U940 ( .A(G2090), .B(G35), .Z(n842) );
  XOR2_X1 U941 ( .A(KEYINPUT54), .B(G34), .Z(n840) );
  XNOR2_X1 U942 ( .A(G2084), .B(n840), .ZN(n841) );
  NAND2_X1 U943 ( .A1(n842), .A2(n841), .ZN(n855) );
  XNOR2_X1 U944 ( .A(G2067), .B(G26), .ZN(n844) );
  XNOR2_X1 U945 ( .A(G33), .B(G2072), .ZN(n843) );
  NOR2_X1 U946 ( .A1(n844), .A2(n843), .ZN(n849) );
  XOR2_X1 U947 ( .A(G1991), .B(G25), .Z(n845) );
  NAND2_X1 U948 ( .A1(n845), .A2(G28), .ZN(n847) );
  XNOR2_X1 U949 ( .A(G32), .B(G1996), .ZN(n846) );
  NOR2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U951 ( .A1(n849), .A2(n848), .ZN(n852) );
  XOR2_X1 U952 ( .A(G27), .B(n850), .Z(n851) );
  NOR2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT53), .ZN(n854) );
  NOR2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n945) );
  XNOR2_X1 U957 ( .A(n856), .B(n945), .ZN(n857) );
  NOR2_X1 U958 ( .A1(G29), .A2(n857), .ZN(n882) );
  XOR2_X1 U959 ( .A(G16), .B(KEYINPUT56), .Z(n858) );
  XNOR2_X1 U960 ( .A(KEYINPUT118), .B(n858), .ZN(n880) );
  XNOR2_X1 U961 ( .A(n1003), .B(G1341), .ZN(n863) );
  XOR2_X1 U962 ( .A(G1966), .B(G168), .Z(n859) );
  NOR2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U964 ( .A(KEYINPUT57), .B(n861), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n874) );
  NAND2_X1 U966 ( .A1(G1971), .A2(G303), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n867) );
  XNOR2_X1 U968 ( .A(G1956), .B(G299), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT119), .B(n872), .Z(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n878) );
  XNOR2_X1 U974 ( .A(n1004), .B(G1348), .ZN(n876) );
  XOR2_X1 U975 ( .A(G301), .B(G1961), .Z(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G11), .A2(n883), .ZN(n912) );
  XOR2_X1 U981 ( .A(G1961), .B(KEYINPUT120), .Z(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(G5), .ZN(n896) );
  XNOR2_X1 U983 ( .A(G1956), .B(G20), .ZN(n886) );
  XNOR2_X1 U984 ( .A(G6), .B(G1981), .ZN(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n893) );
  XOR2_X1 U986 ( .A(KEYINPUT122), .B(G4), .Z(n888) );
  XNOR2_X1 U987 ( .A(G1348), .B(KEYINPUT59), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(KEYINPUT121), .B(n889), .Z(n891) );
  XNOR2_X1 U990 ( .A(G1341), .B(G19), .ZN(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT60), .B(n894), .Z(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n904) );
  XNOR2_X1 U995 ( .A(G1986), .B(G24), .ZN(n898) );
  XNOR2_X1 U996 ( .A(G23), .B(G1976), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n901) );
  XNOR2_X1 U998 ( .A(G1971), .B(KEYINPUT123), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(G22), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(KEYINPUT58), .B(n902), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n906) );
  XOR2_X1 U1003 ( .A(G1966), .B(G21), .Z(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n907), .B(KEYINPUT61), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(KEYINPUT124), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G16), .A2(n909), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT125), .B(n910), .Z(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(KEYINPUT126), .ZN(n949) );
  NAND2_X1 U1011 ( .A1(G139), .A2(n978), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(G103), .A2(n533), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(G127), .A2(n975), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(G115), .A2(n976), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1017 ( .A(KEYINPUT47), .B(n918), .Z(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n989) );
  XOR2_X1 U1019 ( .A(G2072), .B(n989), .Z(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(n921), .ZN(n923) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n924), .Z(n943) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n987), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT113), .B(n930), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT114), .B(n935), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT51), .B(n938), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT115), .B(n941), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT62), .B(n950), .Z(G311) );
  XNOR2_X1 U1043 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(G325) );
  INV_X1 U1045 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1046 ( .A(n953), .B(G2474), .Z(n963) );
  XOR2_X1 U1047 ( .A(KEYINPUT110), .B(G1981), .Z(n955) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G1956), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n955), .B(n954), .ZN(n959) );
  XOR2_X1 U1050 ( .A(KEYINPUT41), .B(G1976), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G1991), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n957), .B(n956), .ZN(n958) );
  XOR2_X1 U1053 ( .A(n959), .B(n958), .Z(n961) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G1971), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n963), .B(n962), .ZN(G229) );
  XNOR2_X1 U1057 ( .A(G2078), .B(G2072), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(G2100), .ZN(n974) );
  XOR2_X1 U1059 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT43), .B(KEYINPUT42), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n966), .B(n965), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT109), .B(G2096), .Z(n968) );
  XNOR2_X1 U1063 ( .A(G2090), .B(G2678), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(n968), .B(n967), .ZN(n969) );
  XOR2_X1 U1065 ( .A(n970), .B(n969), .Z(n972) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G2084), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(G227) );
  NAND2_X1 U1069 ( .A1(G130), .A2(n975), .ZN(n986) );
  NAND2_X1 U1070 ( .A1(n976), .A2(G118), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(KEYINPUT111), .B(n977), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(G142), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(G106), .A2(n533), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1075 ( .A(KEYINPUT112), .B(n981), .Z(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT45), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(n987), .ZN(n999) );
  XNOR2_X1 U1080 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n992), .B(n991), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n993), .B(G162), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G164), .B(G160), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n995), .B(n994), .ZN(n996) );
  XOR2_X1 U1086 ( .A(n997), .B(n996), .Z(n998) );
  XNOR2_X1 U1087 ( .A(n999), .B(n998), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(n1001), .B(n1000), .Z(n1002) );
  NOR2_X1 U1089 ( .A1(G37), .A2(n1002), .ZN(G395) );
  XNOR2_X1 U1090 ( .A(n1003), .B(G286), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(G301), .B(n1004), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(n1008), .B(n1007), .Z(n1009) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1009), .ZN(G397) );
  NAND2_X1 U1095 ( .A1(G319), .A2(n1010), .ZN(n1013) );
  NOR2_X1 U1096 ( .A1(G229), .A2(G227), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(KEYINPUT49), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(G395), .A2(G397), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(G225) );
  INV_X1 U1101 ( .A(G225), .ZN(G308) );
  INV_X1 U1102 ( .A(G57), .ZN(G237) );
  INV_X1 U1103 ( .A(n1016), .ZN(G223) );
endmodule

