//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G71gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G99gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT68), .B1(new_n207), .B2(KEYINPUT27), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(G183gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G183gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT27), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT28), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT27), .B(G183gat), .Z(new_n220));
  OAI21_X1  g019(.A(KEYINPUT28), .B1(new_n220), .B2(G190gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT69), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226));
  OAI22_X1  g025(.A1(new_n226), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n218), .A2(new_n219), .A3(new_n221), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n213), .A2(G183gat), .ZN(new_n233));
  AOI21_X1  g032(.A(G190gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n231), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n225), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT25), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n241), .A2(new_n225), .A3(new_n243), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n222), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT65), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n207), .A2(new_n251), .A3(KEYINPUT64), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n236), .A2(new_n252), .A3(new_n254), .A4(new_n237), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n246), .A2(new_n249), .A3(new_n250), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n230), .A2(new_n245), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G120gat), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(new_n259), .B2(KEYINPUT1), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  INV_X1    g065(.A(G120gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(G113gat), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n263), .B(new_n264), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n260), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT70), .B(new_n261), .C1(new_n259), .C2(KEYINPUT1), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n258), .B1(new_n257), .B2(new_n273), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n230), .A2(new_n272), .A3(new_n245), .A4(new_n256), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT71), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n206), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n204), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n230), .A2(new_n245), .A3(new_n256), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n283), .B2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n274), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n278), .B(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n205), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT73), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n280), .A2(new_n291), .A3(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n280), .B(KEYINPUT32), .C1(new_n281), .C2(new_n204), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(new_n287), .A3(new_n205), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n293), .A2(new_n294), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n293), .B2(new_n294), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(KEYINPUT22), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n315), .B2(KEYINPUT29), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  XNOR2_X1  g116(.A(G141gat), .B(G148gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G155gat), .B(G162gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT2), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n317), .A3(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n331), .A2(new_n317), .A3(new_n322), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n322), .B1(new_n331), .B2(new_n317), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n308), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(KEYINPUT77), .A3(new_n308), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n315), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(G50gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(G50gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT31), .B(G22gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n345), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n345), .B2(new_n346), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n307), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n346), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n349), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n346), .A3(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n306), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G8gat), .B(G36gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G64gat), .ZN(new_n360));
  INV_X1    g159(.A(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n257), .A2(G226gat), .A3(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n257), .A2(new_n365), .B1(G226gat), .B2(G233gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n364), .A2(new_n366), .A3(new_n315), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n257), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n343), .B1(new_n370), .B2(new_n363), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n362), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n315), .B1(new_n364), .B2(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n343), .A3(new_n363), .ZN(new_n374));
  INV_X1    g173(.A(new_n362), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n373), .A2(new_n374), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n377), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT83), .B1(new_n377), .B2(new_n379), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n340), .A2(new_n341), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n272), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n270), .A2(KEYINPUT76), .A3(new_n271), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n334), .A2(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n270), .A2(new_n271), .B1(new_n324), .B2(new_n332), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n272), .A2(new_n333), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n272), .A2(new_n393), .A3(new_n333), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(KEYINPUT79), .A3(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n383), .B(new_n390), .C1(new_n397), .C2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n270), .A2(KEYINPUT76), .A3(new_n271), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT76), .B1(new_n270), .B2(new_n271), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n395), .B1(new_n407), .B2(new_n333), .ZN(new_n408));
  INV_X1    g207(.A(new_n383), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT0), .B(G57gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  AOI22_X1  g214(.A1(new_n386), .A2(new_n387), .B1(new_n334), .B2(KEYINPUT3), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n416), .A2(new_n384), .B1(new_n398), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n418), .A2(new_n404), .A3(new_n383), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n411), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT80), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n411), .A2(new_n419), .ZN(new_n422));
  INV_X1    g221(.A(new_n415), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n411), .A2(new_n426), .A3(new_n415), .A4(new_n419), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n424), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n415), .B1(new_n411), .B2(new_n419), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT35), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n305), .A2(new_n358), .A3(new_n382), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n430), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n377), .A2(new_n379), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI211_X1 g236(.A(KEYINPUT81), .B(new_n435), .C1(new_n428), .C2(new_n430), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n358), .B1(new_n302), .B2(new_n303), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT35), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT37), .B1(new_n367), .B2(new_n371), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT37), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n373), .A2(new_n374), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n362), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n445), .B2(KEYINPUT84), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n376), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n428), .A2(new_n430), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n383), .B(new_n395), .C1(new_n407), .C2(new_n333), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(KEYINPUT39), .C1(new_n418), .C2(new_n383), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n418), .A2(new_n383), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n415), .C1(new_n456), .C2(KEYINPUT39), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n429), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n457), .A2(new_n453), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n458), .B(new_n459), .C1(new_n380), .C2(new_n381), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n452), .A2(new_n460), .A3(new_n358), .ZN(new_n461));
  INV_X1    g260(.A(new_n303), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n293), .A2(new_n301), .A3(new_n294), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n302), .B2(new_n303), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n358), .B(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n437), .B2(new_n438), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n442), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G57gat), .B(G64gat), .Z(new_n474));
  INV_X1    g273(.A(KEYINPUT9), .ZN(new_n475));
  INV_X1    g274(.A(G71gat), .ZN(new_n476));
  INV_X1    g275(.A(G78gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G78gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n480), .B(KEYINPUT91), .Z(new_n481));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n479), .B(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n474), .A2(new_n478), .ZN(new_n484));
  OR3_X1    g283(.A1(new_n483), .A2(KEYINPUT90), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT90), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n487), .A2(KEYINPUT21), .ZN(new_n488));
  XOR2_X1   g287(.A(G127gat), .B(G155gat), .Z(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(KEYINPUT21), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT16), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(G1gat), .B2(new_n492), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(G8gat), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n501));
  INV_X1    g300(.A(G231gat), .ZN(new_n502));
  INV_X1    g301(.A(G233gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n500), .B2(new_n501), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n490), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n507), .ZN(new_n509));
  INV_X1    g308(.A(new_n490), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n513));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n511), .A3(new_n515), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n521), .B(new_n523), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  XOR2_X1   g323(.A(G43gat), .B(G50gat), .Z(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(KEYINPUT86), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT7), .B1(new_n534), .B2(KEYINPUT93), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT95), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n537), .B(KEYINPUT7), .C1(new_n534), .C2(KEYINPUT93), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT93), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT96), .B(G92gat), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n543), .A2(new_n544), .B1(KEYINPUT8), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n536), .A2(KEYINPUT93), .A3(new_n540), .A4(new_n538), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G99gat), .B(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n542), .A2(new_n549), .A3(new_n546), .A4(new_n547), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT41), .ZN(new_n558));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .C1(new_n556), .C2(new_n530), .ZN(new_n560));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n558), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n561), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n560), .B(new_n561), .ZN(new_n568));
  INV_X1    g367(.A(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n517), .A2(new_n518), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n473), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G204gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT101), .ZN(new_n575));
  INV_X1    g374(.A(G176gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT10), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n549), .B(KEYINPUT99), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n548), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n487), .B(new_n583), .C1(new_n554), .C2(new_n555), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n485), .A2(new_n486), .ZN(new_n585));
  INV_X1    g384(.A(new_n481), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n556), .A2(KEYINPUT98), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT98), .B1(new_n556), .B2(new_n587), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n581), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  OR3_X1    g389(.A1(new_n556), .A2(new_n587), .A3(new_n581), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n580), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n556), .A2(new_n587), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n587), .A3(KEYINPUT98), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(new_n579), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n592), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n578), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n598), .A2(new_n579), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n590), .A2(new_n591), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n605), .B(KEYINPUT100), .C1(new_n606), .C2(new_n580), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(new_n577), .A3(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n497), .A2(new_n530), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n497), .A2(new_n530), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  AOI211_X1 g416(.A(KEYINPUT87), .B(new_n615), .C1(new_n611), .C2(new_n612), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n531), .A2(new_n497), .A3(new_n532), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n614), .A4(new_n611), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n614), .A3(new_n611), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n619), .A2(new_n621), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n621), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n635), .A3(KEYINPUT88), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT88), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n637), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n609), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n572), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n434), .B(KEYINPUT102), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n493), .ZN(G1324gat));
  INV_X1    g444(.A(new_n641), .ZN(new_n646));
  INV_X1    g445(.A(new_n382), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n649));
  AND2_X1   g448(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(G8gat), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT42), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(G1325gat));
  AOI21_X1  g455(.A(G15gat), .B1(new_n646), .B2(new_n305), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n464), .A2(new_n466), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(G15gat), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n358), .A2(new_n469), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT82), .B1(new_n353), .B2(new_n357), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n570), .A2(new_n567), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n442), .B2(new_n472), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n517), .A2(new_n518), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n640), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n519), .A3(new_n642), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n473), .B2(new_n668), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n434), .A2(new_n436), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT81), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n434), .A2(new_n433), .A3(new_n436), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n663), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT105), .B1(new_n679), .B2(new_n467), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n471), .A2(new_n681), .A3(new_n658), .A4(new_n461), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n442), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n667), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n609), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT104), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n639), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n670), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n643), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n693), .ZN(G1328gat));
  NOR3_X1   g493(.A1(new_n671), .A2(G36gat), .A3(new_n382), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n692), .B2(new_n382), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n692), .B2(new_n658), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n671), .A2(G43gat), .A3(new_n304), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT47), .B1(new_n700), .B2(KEYINPUT107), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1330gat));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(G50gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n692), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n470), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n672), .A2(new_n705), .A3(new_n470), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n358), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n686), .A2(new_n670), .A3(new_n711), .A4(new_n691), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(new_n708), .ZN(new_n714));
  OAI221_X1 g513(.A(new_n704), .B1(new_n707), .B2(new_n710), .C1(new_n714), .C2(new_n709), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n707), .A2(new_n710), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n709), .B1(new_n713), .B2(new_n708), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n639), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n571), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n683), .A2(new_n690), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n642), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n647), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT49), .B(G64gat), .Z(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(G1333gat));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n476), .A3(new_n305), .ZN(new_n729));
  INV_X1    g528(.A(new_n658), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n476), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n470), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  INV_X1    g535(.A(new_n670), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n720), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n609), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n675), .B2(new_n685), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741), .B2(new_n643), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n683), .A2(new_n667), .A3(new_n738), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n683), .A2(KEYINPUT51), .A3(new_n667), .A4(new_n738), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n747), .A2(new_n746), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n609), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n642), .A2(new_n544), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n742), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n747), .ZN(new_n753));
  INV_X1    g552(.A(new_n690), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(G92gat), .A3(new_n382), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n543), .B1(new_n740), .B2(new_n647), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT52), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n748), .A2(new_n749), .A3(new_n755), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n741), .B2(new_n658), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n304), .A2(G99gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n750), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT111), .ZN(G1338gat));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  INV_X1    g566(.A(G106gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n690), .A2(new_n768), .A3(new_n711), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n753), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g570(.A(KEYINPUT112), .B(new_n769), .C1(new_n745), .C2(new_n747), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n768), .B1(new_n740), .B2(new_n470), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n766), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G106gat), .B1(new_n741), .B2(new_n358), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n748), .A2(new_n749), .A3(new_n770), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n766), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT113), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n778), .A3(new_n766), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n774), .A2(new_n771), .A3(new_n772), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n782), .C1(new_n783), .C2(new_n766), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n784), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n578), .B1(new_n592), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n590), .A2(new_n580), .A3(new_n591), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n592), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n787), .B(KEYINPUT55), .C1(new_n592), .C2(new_n789), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n792), .A2(new_n720), .A3(new_n604), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n614), .B1(new_n620), .B2(new_n611), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n613), .A2(new_n616), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n629), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n631), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n609), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n667), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n604), .A2(new_n793), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n798), .B1(new_n570), .B2(new_n567), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(new_n792), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n670), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n571), .A2(new_n609), .A3(new_n720), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n470), .A2(new_n647), .A3(new_n304), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n642), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n639), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n802), .A2(new_n792), .A3(new_n803), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n639), .B1(new_n791), .B2(new_n790), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n802), .A2(new_n813), .B1(new_n609), .B2(new_n799), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n667), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n806), .B1(new_n815), .B2(new_n670), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n643), .A3(new_n439), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n382), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n720), .A2(new_n265), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n811), .B1(new_n818), .B2(new_n819), .ZN(G1340gat));
  INV_X1    g619(.A(new_n818), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n267), .A3(new_n609), .ZN(new_n822));
  OAI21_X1  g621(.A(G120gat), .B1(new_n810), .B2(new_n754), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n825), .A3(new_n670), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n821), .A2(KEYINPUT114), .A3(new_n737), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT114), .B1(new_n821), .B2(new_n737), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n829), .B2(new_n825), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n817), .A2(new_n831), .A3(new_n667), .A4(new_n382), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT56), .Z(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n810), .B2(new_n668), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1343gat));
  AOI21_X1  g634(.A(new_n358), .B1(new_n805), .B2(new_n807), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(new_n839), .C1(new_n816), .C2(new_n358), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n790), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n720), .A3(new_n604), .A4(new_n793), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n667), .B1(new_n843), .B2(new_n800), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n804), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n807), .B1(new_n845), .B2(new_n737), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT57), .A3(new_n470), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n837), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n730), .A2(new_n643), .A3(new_n647), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(G141gat), .A3(new_n720), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n816), .A2(new_n643), .A3(new_n358), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n730), .A2(new_n647), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n327), .B1(new_n854), .B2(new_n639), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n851), .A2(KEYINPUT58), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1344gat));
  NOR3_X1   g659(.A1(new_n854), .A2(G148gat), .A3(new_n687), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n844), .B2(new_n804), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n639), .B1(new_n790), .B2(new_n841), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n802), .A2(new_n865), .B1(new_n609), .B2(new_n799), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n864), .B(new_n812), .C1(new_n866), .C2(new_n667), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n867), .A3(new_n670), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n806), .B(KEYINPUT117), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n663), .A2(KEYINPUT57), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n808), .A2(new_n711), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n872), .A2(new_n874), .A3(new_n609), .A4(new_n849), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G148gat), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT59), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n848), .A2(new_n609), .A3(new_n849), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n328), .A2(KEYINPUT59), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT119), .B(new_n862), .C1(new_n877), .C2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n876), .A2(KEYINPUT59), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n861), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1345gat));
  INV_X1    g684(.A(new_n854), .ZN(new_n886));
  AOI21_X1  g685(.A(G155gat), .B1(new_n886), .B2(new_n737), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n737), .A2(G155gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n850), .B2(new_n888), .ZN(G1346gat));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n667), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G162gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n668), .A2(G162gat), .A3(new_n647), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n852), .A2(new_n658), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT120), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n642), .A2(new_n382), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n816), .A2(new_n439), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(G169gat), .A3(new_n639), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n816), .A2(new_n897), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n663), .A3(new_n305), .ZN(new_n903));
  OAI21_X1  g702(.A(G169gat), .B1(new_n903), .B2(new_n639), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n898), .B2(new_n609), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n903), .A2(new_n576), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n690), .ZN(G1349gat));
  NOR2_X1   g707(.A1(new_n214), .A2(new_n215), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n903), .B2(new_n670), .ZN(new_n910));
  INV_X1    g709(.A(new_n220), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n898), .A2(new_n737), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n914), .A2(KEYINPUT60), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT60), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n903), .B2(new_n668), .ZN(new_n920));
  XOR2_X1   g719(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n251), .A3(new_n667), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  NAND4_X1  g723(.A1(new_n872), .A2(new_n874), .A3(new_n658), .A4(new_n896), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n925), .A2(KEYINPUT124), .A3(new_n639), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT124), .B1(new_n925), .B2(new_n639), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(G197gat), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n896), .A2(new_n658), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n873), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G197gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n720), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(G1352gat));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(G204gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n609), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  NOR2_X1   g735(.A1(new_n925), .A2(new_n754), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n934), .ZN(G1353gat));
  NAND3_X1  g737(.A1(new_n930), .A2(new_n310), .A3(new_n737), .ZN(new_n939));
  INV_X1    g738(.A(new_n871), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n868), .B2(new_n869), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n836), .A2(new_n839), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(new_n929), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n737), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n939), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  AOI21_X1  g746(.A(new_n668), .B1(new_n943), .B2(KEYINPUT126), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n925), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n311), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n311), .A3(new_n667), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n667), .B1(new_n925), .B2(new_n949), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n943), .A2(KEYINPUT126), .ZN(new_n956));
  OAI21_X1  g755(.A(G218gat), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n958), .A3(new_n952), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n954), .A2(new_n959), .ZN(G1355gat));
endmodule


