//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT75), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT81), .B(G155gat), .Z(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G162gat), .ZN(new_n223));
  XOR2_X1   g022(.A(G141gat), .B(G148gat), .Z(new_n224));
  XNOR2_X1  g023(.A(G155gat), .B(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(KEYINPUT80), .ZN(new_n229));
  NOR2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n228), .B(new_n229), .C1(KEYINPUT80), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n219), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n232), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(G228gat), .A3(G233gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G228gat), .A2(G233gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n210), .A2(new_n211), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n213), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT3), .B1(new_n245), .B2(new_n234), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n236), .B(new_n243), .C1(new_n240), .C2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT31), .B(G50gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n242), .B2(new_n247), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n204), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n203), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n257));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT65), .Z(new_n259));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n260), .A2(KEYINPUT23), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(KEYINPUT23), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n257), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n260), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT23), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n261), .A2(KEYINPUT25), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n268), .A4(new_n259), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n259), .A2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(G183gat), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n288), .A2(KEYINPUT27), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n283), .B(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G190gat), .ZN(new_n293));
  OAI221_X1 g092(.A(new_n265), .B1(new_n285), .B2(new_n290), .C1(new_n293), .C2(new_n286), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n276), .B1(new_n282), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G226gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n295), .B2(new_n234), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n220), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n293), .A2(new_n286), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n265), .B1(new_n290), .B2(new_n285), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n279), .A2(new_n281), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n305), .A2(new_n306), .B1(new_n270), .B2(new_n275), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT29), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n299), .B(new_n237), .C1(new_n308), .C2(new_n298), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT37), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n302), .A2(new_n309), .A3(KEYINPUT86), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n298), .B1(new_n295), .B2(new_n238), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n316), .A3(new_n220), .ZN(new_n317));
  INV_X1    g116(.A(new_n234), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n307), .A2(new_n318), .B1(new_n296), .B2(new_n297), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n237), .B1(new_n319), .B2(new_n299), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT77), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n309), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(KEYINPUT37), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n315), .A2(new_n324), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT38), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n327), .B(KEYINPUT78), .Z(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(KEYINPUT38), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n237), .B1(new_n300), .B2(new_n301), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT37), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n300), .A2(new_n316), .A3(new_n237), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n313), .B2(new_n314), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  OR3_X1    g142(.A1(new_n343), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT70), .B1(new_n343), .B2(G113gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(G120gat), .ZN(new_n347));
  XOR2_X1   g146(.A(G127gat), .B(G134gat), .Z(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT1), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n346), .A2(G120gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n343), .A2(G113gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n353), .B2(KEYINPUT1), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n232), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT82), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(new_n232), .B2(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n232), .A2(new_n355), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n342), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n355), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n233), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(new_n359), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(KEYINPUT4), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n367), .A2(new_n342), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(new_n369), .B2(KEYINPUT4), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n341), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT6), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n302), .A2(new_n309), .A3(new_n327), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n375), .ZN(new_n380));
  INV_X1    g179(.A(new_n341), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n377), .B(new_n378), .C1(new_n382), .C2(new_n376), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n337), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n256), .B1(new_n330), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n331), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n321), .A2(new_n323), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT30), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n378), .A2(new_n390), .A3(new_n388), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n378), .B2(new_n388), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n387), .B(new_n389), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT40), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n233), .A2(new_n366), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n362), .B1(new_n374), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n361), .B2(new_n363), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n341), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT39), .B(new_n362), .C1(new_n374), .C2(new_n395), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT84), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n376), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT84), .B1(new_n398), .B2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT40), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n393), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n393), .A2(new_n402), .A3(KEYINPUT85), .A4(new_n404), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT71), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n307), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n355), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n295), .A2(KEYINPUT71), .A3(new_n365), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(G227gat), .A3(G233gat), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n412), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(KEYINPUT32), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n418), .B(KEYINPUT32), .C1(new_n419), .C2(new_n412), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n417), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT34), .ZN(new_n426));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n426), .B1(new_n425), .B2(new_n427), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n422), .A3(new_n423), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n424), .B2(new_n431), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n430), .A2(new_n422), .A3(new_n423), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n430), .B1(new_n423), .B2(new_n422), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n436), .B(new_n439), .C1(new_n442), .C2(KEYINPUT72), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n376), .B1(new_n382), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT83), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n377), .ZN(new_n448));
  INV_X1    g247(.A(new_n393), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n256), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n409), .A2(new_n435), .A3(new_n443), .A4(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n253), .A2(new_n255), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n432), .A3(new_n433), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT35), .B1(new_n454), .B2(new_n450), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n438), .B1(new_n434), .B2(new_n437), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  MUX2_X1   g256(.A(new_n382), .B(new_n379), .S(new_n376), .Z(new_n458));
  NOR3_X1   g257(.A1(new_n256), .A2(new_n458), .A3(KEYINPUT35), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n449), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(G36gat), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n466));
  OAI21_X1  g265(.A(G29gat), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n468), .B(new_n469), .C1(G29gat), .C2(G36gat), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT91), .B(KEYINPUT15), .ZN(new_n472));
  OR2_X1    g271(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n474));
  AOI21_X1  g273(.A(G50gat), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G50gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT93), .B1(new_n476), .B2(G43gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n478));
  INV_X1    g277(.A(G43gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n479), .A3(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n472), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(G43gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(G50gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT15), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n465), .A3(KEYINPUT88), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n468), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT14), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n471), .A2(new_n482), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n467), .A2(new_n489), .A3(new_n470), .ZN(new_n491));
  INV_X1    g290(.A(new_n485), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n491), .A2(KEYINPUT90), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT90), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n490), .B(KEYINPUT17), .C1(new_n493), .C2(new_n494), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(G1gat), .ZN(new_n501));
  INV_X1    g300(.A(G15gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G22gat), .ZN(new_n503));
  INV_X1    g302(.A(G22gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G15gat), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G1gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n503), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT95), .A3(new_n499), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT94), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n514), .B2(new_n499), .ZN(new_n518));
  INV_X1    g317(.A(new_n508), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT94), .A3(G8gat), .A4(new_n512), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n516), .B2(new_n521), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n497), .B(new_n498), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT97), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n516), .A2(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT96), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n498), .A4(new_n497), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n495), .A2(new_n527), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT98), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT99), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n538), .B1(new_n526), .B2(new_n532), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(KEYINPUT18), .ZN(new_n545));
  INV_X1    g344(.A(new_n534), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n495), .A2(new_n527), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n536), .B(KEYINPUT13), .Z(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n544), .B2(KEYINPUT18), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT11), .B(G169gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n545), .A3(new_n551), .A4(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n539), .ZN(new_n560));
  INV_X1    g359(.A(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n544), .A2(KEYINPUT18), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n497), .A2(new_n498), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  INV_X1    g369(.A(G92gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G99gat), .B(G106gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n495), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT104), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT103), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G57gat), .A2(G64gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT101), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT101), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n603), .A2(new_n604), .B1(KEYINPUT9), .B2(new_n595), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n592), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n591), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT102), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n596), .B1(new_n613), .B2(new_n602), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n614), .A2(new_n615), .A3(new_n609), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n599), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(G127gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n620), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n619), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G127gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n527), .B1(new_n618), .B2(KEYINPUT21), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n622), .B2(new_n626), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n629), .B2(new_n631), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n588), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n297), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n617), .A2(new_n576), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n605), .A2(KEYINPUT102), .A3(new_n610), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n615), .B1(new_n614), .B2(new_n609), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n599), .A3(new_n575), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n647), .A2(new_n599), .A3(new_n575), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT10), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n642), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n642), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n643), .B2(new_n648), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n652), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n652), .B2(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AND4_X1   g461(.A1(new_n462), .A2(new_n565), .A3(new_n640), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n448), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n663), .A2(new_n393), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n499), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(G1325gat));
  NAND3_X1  g472(.A1(new_n663), .A2(new_n502), .A3(new_n456), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n443), .A2(new_n435), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n663), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n676), .B2(new_n502), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n256), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n588), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n452), .B2(new_n461), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n637), .A2(new_n639), .ZN(new_n683));
  INV_X1    g482(.A(new_n565), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(new_n684), .A3(new_n661), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n486), .A3(new_n664), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n462), .A2(new_n588), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n685), .B(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n448), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n689), .A2(new_n697), .ZN(G1328gat));
  NOR4_X1   g497(.A1(new_n686), .A2(new_n449), .A3(new_n464), .A4(new_n466), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n696), .A2(new_n449), .B1(new_n464), .B2(new_n466), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1329gat));
  OAI211_X1 g501(.A(new_n473), .B(new_n474), .C1(new_n686), .C2(new_n457), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n473), .A2(new_n474), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n675), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT47), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n708), .B(new_n703), .C1(new_n696), .C2(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1330gat));
  NAND4_X1  g509(.A1(new_n692), .A2(new_n256), .A3(new_n693), .A4(new_n695), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G50gat), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT48), .B1(new_n712), .B2(KEYINPUT106), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n687), .A2(new_n476), .A3(new_n256), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n712), .B(new_n714), .C1(KEYINPUT106), .C2(KEYINPUT48), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  AND4_X1   g517(.A1(new_n462), .A2(new_n684), .A3(new_n640), .A4(new_n661), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n664), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n393), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT49), .B(G64gat), .Z(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n722), .B2(new_n724), .ZN(G1333gat));
  AOI21_X1  g524(.A(new_n589), .B1(new_n719), .B2(new_n675), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n457), .A2(G71gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n719), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n719), .A2(new_n256), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n683), .A2(new_n565), .A3(new_n662), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n694), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n448), .ZN(new_n734));
  NAND2_X1  g533(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n683), .A2(new_n565), .A3(new_n736), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n462), .A2(new_n588), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n682), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n664), .A2(new_n570), .A3(new_n661), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  NAND4_X1  g542(.A1(new_n692), .A2(new_n393), .A3(new_n693), .A4(new_n732), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n449), .A2(G92gat), .A3(new_n662), .ZN(new_n745));
  AOI22_X1  g544(.A1(G92gat), .A2(new_n744), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT108), .B1(new_n744), .B2(G92gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT52), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(G92gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n740), .A2(new_n745), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(KEYINPUT52), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n748), .A2(new_n753), .ZN(G1337gat));
  INV_X1    g553(.A(new_n675), .ZN(new_n755));
  OAI21_X1  g554(.A(G99gat), .B1(new_n733), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n457), .A2(G99gat), .A3(new_n662), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT109), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n741), .B2(new_n758), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n692), .A2(new_n256), .A3(new_n693), .A4(new_n732), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n453), .A2(G106gat), .A3(new_n662), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n740), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT53), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n761), .B(new_n763), .C1(KEYINPUT110), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1339gat));
  AND3_X1   g568(.A1(new_n640), .A2(new_n684), .A3(new_n662), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n575), .B1(new_n647), .B2(new_n599), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n650), .A2(new_n772), .A3(KEYINPUT10), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n648), .A2(new_n644), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n653), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n649), .A2(new_n651), .A3(new_n642), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n657), .B1(new_n652), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(KEYINPUT55), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n659), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT55), .B1(new_n777), .B2(new_n779), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n531), .B1(new_n566), .B2(new_n530), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n525), .A2(KEYINPUT97), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n534), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(new_n787), .A3(new_n536), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n548), .A2(new_n549), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n546), .B1(new_n526), .B2(new_n532), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT111), .B1(new_n790), .B2(new_n537), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n555), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n588), .A2(new_n783), .A3(new_n558), .A4(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT99), .B1(new_n540), .B2(new_n541), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n544), .A2(new_n543), .A3(KEYINPUT18), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n562), .A2(new_n559), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n662), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n793), .B1(new_n565), .B2(new_n783), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n588), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n565), .A2(new_n783), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n558), .A3(new_n661), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT112), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n795), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n771), .B1(new_n808), .B2(new_n683), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n448), .A2(new_n393), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n453), .A2(new_n809), .A3(new_n456), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n346), .B1(new_n811), .B2(new_n565), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT113), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n804), .A2(new_n805), .A3(new_n802), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n681), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n794), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n683), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n770), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n448), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n454), .A2(new_n393), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n565), .A2(new_n346), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n661), .A3(new_n821), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n662), .A2(new_n343), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n343), .A2(new_n825), .B1(new_n811), .B2(new_n826), .ZN(G1341gat));
  AOI21_X1  g626(.A(new_n625), .B1(new_n811), .B2(new_n683), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n822), .A2(G127gat), .A3(new_n818), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n828), .A2(new_n829), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n811), .B2(new_n588), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT114), .Z(new_n833));
  NOR3_X1   g632(.A1(new_n822), .A2(G134gat), .A3(new_n681), .ZN(new_n834));
  NAND2_X1  g633(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n837));
  OAI211_X1 g636(.A(new_n833), .B(new_n836), .C1(new_n834), .C2(new_n837), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n755), .A2(new_n810), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n794), .B1(new_n801), .B2(new_n588), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n818), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n770), .B1(new_n841), .B2(KEYINPUT116), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(KEYINPUT116), .B2(new_n841), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n453), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n819), .B2(new_n453), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(G141gat), .A3(new_n565), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n755), .B2(new_n256), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n675), .A2(KEYINPUT117), .A3(new_n453), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n393), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n820), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n684), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n849), .B1(new_n855), .B2(G141gat), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n856), .B(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(new_n854), .ZN(new_n859));
  INV_X1    g658(.A(G148gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n661), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n453), .B1(new_n771), .B2(new_n841), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n863), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n809), .A2(new_n845), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n867), .A2(new_n755), .A3(new_n661), .A4(new_n810), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n862), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT59), .B(new_n860), .C1(new_n848), .C2(new_n661), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n861), .B1(new_n869), .B2(new_n870), .ZN(G1345gat));
  INV_X1    g670(.A(new_n222), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n859), .A2(new_n872), .A3(new_n683), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n848), .A2(new_n683), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n872), .ZN(G1346gat));
  AOI21_X1  g674(.A(G162gat), .B1(new_n859), .B2(new_n588), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n588), .A2(G162gat), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n876), .B1(new_n848), .B2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n454), .A2(new_n449), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT120), .Z(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n819), .B2(new_n664), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n807), .A2(new_n681), .A3(new_n814), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n683), .B1(new_n883), .B2(new_n794), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n448), .C1(new_n884), .C2(new_n770), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n565), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n819), .A2(new_n256), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n664), .A2(new_n449), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n457), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n565), .A2(G169gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(G1348gat));
  INV_X1    g693(.A(G176gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n895), .A3(new_n661), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n892), .A2(new_n661), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n895), .ZN(G1349gat));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n809), .A2(new_n453), .A3(new_n683), .A4(new_n891), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT121), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n888), .A2(new_n902), .A3(new_n683), .A4(new_n891), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n903), .A3(G183gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n818), .A2(new_n292), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT122), .A3(KEYINPUT123), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n288), .B1(new_n900), .B2(KEYINPUT121), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n903), .A2(new_n910), .B1(new_n886), .B2(new_n905), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT60), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n899), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n904), .A2(new_n906), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n907), .B1(new_n917), .B2(KEYINPUT123), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(KEYINPUT124), .A3(new_n909), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1350gat));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n892), .A2(new_n588), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(G190gat), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT61), .B(new_n287), .C1(new_n892), .C2(new_n588), .ZN(new_n925));
  INV_X1    g724(.A(new_n886), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n588), .A2(new_n287), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n924), .A2(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI221_X1 g729(.A(KEYINPUT125), .B1(new_n926), .B2(new_n927), .C1(new_n924), .C2(new_n925), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n675), .A2(new_n890), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n867), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n684), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n882), .A2(new_n885), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n675), .A2(new_n449), .A3(new_n453), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n565), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n935), .A2(new_n941), .ZN(G1352gat));
  XOR2_X1   g741(.A(KEYINPUT126), .B(G204gat), .Z(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n662), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n867), .A2(new_n661), .A3(new_n933), .ZN(new_n947));
  AOI22_X1  g746(.A1(new_n946), .A2(KEYINPUT62), .B1(new_n947), .B2(new_n944), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  INV_X1    g748(.A(new_n946), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n946), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n207), .A3(new_n683), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n867), .A2(new_n683), .A3(new_n933), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n934), .B2(new_n681), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n939), .A2(new_n208), .A3(new_n588), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


