//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT0), .B(G128), .Z(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(G146), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G143), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n199), .A2(KEYINPUT65), .A3(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n188), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT11), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G134), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n205), .B2(G134), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n202), .A3(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n203), .A2(new_n206), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n208), .A4(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n192), .A2(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n199), .B2(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT0), .A3(G128), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n201), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(new_n205), .B2(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n205), .A2(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n205), .A2(KEYINPUT67), .A3(G134), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n227));
  OAI21_X1  g041(.A(G128), .B1(new_n227), .B2(new_n217), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n198), .B2(new_n200), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(G128), .A3(new_n227), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G116), .B(G119), .Z(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n220), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT30), .B1(new_n220), .B2(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(new_n226), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n239));
  INV_X1    g053(.A(new_n217), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n194), .A2(G143), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n189), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n190), .B1(new_n244), .B2(KEYINPUT65), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n196), .A2(new_n197), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n193), .A2(new_n195), .A3(G146), .ZN(new_n248));
  AND4_X1   g062(.A1(G128), .A2(new_n248), .A3(new_n240), .A4(new_n227), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n237), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n201), .A2(new_n216), .A3(new_n219), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n236), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n235), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G210), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n258), .B(KEYINPUT27), .Z(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT31), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n220), .A2(new_n231), .A3(KEYINPUT30), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n234), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n235), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n262), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n255), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n235), .A2(KEYINPUT28), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n234), .B1(new_n220), .B2(new_n231), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(new_n262), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT32), .B(new_n187), .C1(new_n273), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n278), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n270), .B2(new_n271), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n284), .B2(new_n263), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT69), .B1(new_n255), .B2(new_n262), .ZN(new_n288));
  AND4_X1   g102(.A1(KEYINPUT69), .A2(new_n266), .A3(new_n267), .A4(new_n262), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT31), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n263), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n187), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(new_n277), .B2(new_n262), .ZN(new_n296));
  INV_X1    g110(.A(new_n255), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n261), .ZN(new_n298));
  AOI21_X1  g112(.A(G902), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n276), .A2(new_n300), .A3(KEYINPUT28), .ZN(new_n301));
  INV_X1    g115(.A(new_n274), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n295), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n281), .A2(new_n286), .A3(new_n294), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT72), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n285), .A2(new_n187), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(new_n287), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n281), .A4(new_n286), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G217), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(G234), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(KEYINPUT16), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n189), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n320), .B(G146), .C1(KEYINPUT16), .C2(new_n322), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n238), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(new_n330), .C1(G119), .C2(new_n238), .ZN(new_n331));
  XNOR2_X1  g145(.A(G119), .B(G128), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT24), .B(G110), .Z(new_n333));
  AOI22_X1  g147(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT73), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n319), .A2(new_n189), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n325), .A3(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT22), .B(G137), .Z(new_n340));
  AND3_X1   g154(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n336), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n336), .B2(new_n339), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n317), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT25), .B1(new_n345), .B2(new_n317), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n318), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n318), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n353));
  INV_X1    g167(.A(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(G104), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT75), .A3(G107), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n354), .A2(KEYINPUT3), .A3(G104), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT3), .B1(new_n354), .B2(G104), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n355), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n356), .B2(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n354), .A2(KEYINPUT3), .A3(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n355), .A4(new_n357), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n369), .A3(G101), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n234), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(KEYINPUT5), .A3(G119), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT82), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n375), .B(G113), .C1(new_n376), .C2(new_n232), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n356), .A2(G107), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n354), .A2(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n367), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n232), .A2(new_n233), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G122), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n372), .A2(new_n384), .A3(new_n386), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n229), .A2(new_n321), .A3(new_n230), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n201), .A2(new_n219), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n321), .ZN(new_n395));
  INV_X1    g209(.A(G224), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G953), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n395), .B(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT7), .B1(new_n396), .B2(G953), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n377), .A2(new_n383), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n381), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n384), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n386), .B(KEYINPUT8), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n400), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n401), .A2(new_n389), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n317), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n399), .A2(new_n317), .A3(new_n410), .A4(new_n408), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(KEYINPUT83), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT81), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n256), .A2(new_n257), .A3(G143), .A4(G214), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n193), .A2(new_n195), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G131), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT86), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n326), .B1(new_n425), .B2(KEYINPUT17), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n424), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT17), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n423), .A2(G131), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n356), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n435), .B(new_n214), .C1(new_n423), .C2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n423), .A2(KEYINPUT85), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n319), .B(new_n189), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n435), .B2(new_n214), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n432), .A2(new_n434), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n434), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n319), .B(KEYINPUT19), .Z(new_n447));
  OAI21_X1  g261(.A(new_n325), .B1(new_n447), .B2(G146), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n428), .B2(new_n430), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT20), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n444), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n434), .B1(new_n432), .B2(new_n443), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n317), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n257), .A2(G952), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(G234), .B2(G237), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n317), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(G898), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n238), .A2(G143), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n421), .B2(new_n238), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G134), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n373), .A2(G122), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n354), .B1(new_n472), .B2(KEYINPUT14), .ZN(new_n473));
  XNOR2_X1  g287(.A(G116), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n199), .A2(new_n477), .A3(G128), .ZN(new_n478));
  OAI211_X1 g292(.A(G134), .B(new_n478), .C1(new_n470), .C2(new_n477), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT87), .B(G107), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n474), .B(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n479), .B(new_n481), .C1(G134), .C2(new_n470), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n316), .A3(G953), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n476), .A2(new_n482), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n317), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n490), .A2(new_n496), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n462), .A2(new_n468), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n352), .A2(new_n419), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G221), .ZN(new_n502));
  INV_X1    g316(.A(new_n484), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n317), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G469), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT76), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n238), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n218), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n248), .A2(new_n240), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT1), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n421), .B2(new_n189), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT76), .B(new_n510), .C1(new_n512), .C2(new_n238), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n230), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT10), .B1(new_n514), .B2(new_n382), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n367), .A2(KEYINPUT10), .A3(new_n380), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n247), .B2(new_n249), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n368), .A2(new_n201), .A3(new_n219), .A4(new_n370), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n216), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n510), .B1(new_n512), .B2(new_n238), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n249), .B1(new_n526), .B2(new_n507), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n381), .B1(new_n527), .B2(new_n513), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n247), .A2(new_n382), .A3(new_n249), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n523), .A2(new_n524), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n521), .A2(new_n522), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT78), .ZN(new_n533));
  OAI221_X1 g347(.A(new_n525), .B1(new_n523), .B2(new_n524), .C1(new_n528), .C2(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n537), .A2(G128), .B1(new_n240), .B2(new_n248), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n230), .B1(new_n538), .B2(KEYINPUT76), .ZN(new_n539));
  INV_X1    g353(.A(new_n513), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n382), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n516), .B1(new_n229), .B2(new_n230), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n371), .B2(new_n394), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n522), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n546), .A3(new_n534), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G110), .B(G140), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n257), .A2(G227), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT74), .Z(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT79), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n216), .B1(new_n515), .B2(new_n520), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT79), .B(new_n216), .C1(new_n515), .C2(new_n520), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n506), .B1(new_n561), .B2(new_n317), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n563));
  INV_X1    g377(.A(new_n553), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n535), .B2(new_n548), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n559), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT80), .B(G469), .C1(new_n566), .C2(G902), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n557), .A2(new_n552), .A3(new_n558), .ZN(new_n568));
  INV_X1    g382(.A(new_n552), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n536), .A2(new_n546), .A3(new_n534), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n506), .A3(new_n317), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n505), .B1(new_n563), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n315), .A2(new_n501), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  OAI21_X1  g391(.A(G472), .B1(new_n292), .B2(G902), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT89), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n295), .B1(new_n285), .B2(new_n317), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n311), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR4_X1   g396(.A1(new_n574), .A2(new_n352), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT33), .B1(new_n485), .B2(KEYINPUT90), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n489), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n489), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n491), .ZN(new_n589));
  NAND2_X1  g403(.A1(G478), .A2(G902), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n490), .B2(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n457), .A2(new_n461), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n468), .ZN(new_n594));
  INV_X1    g408(.A(new_n416), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n412), .B2(new_n413), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n583), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n356), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  OR2_X1    g416(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n603));
  INV_X1    g417(.A(new_n499), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n603), .A2(new_n461), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n467), .B(KEYINPUT93), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n583), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n582), .A2(new_n579), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n336), .A2(new_n339), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT36), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n342), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n614), .B(new_n616), .Z(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n349), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n348), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n620), .A2(new_n500), .A3(new_n419), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n575), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT94), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  AOI21_X1  g439(.A(new_n574), .B1(new_n310), .B2(new_n314), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n596), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT95), .B(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n464), .B1(new_n465), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n606), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  XOR2_X1   g446(.A(new_n629), .B(KEYINPUT39), .Z(new_n633));
  NAND2_X1  g447(.A1(new_n575), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n281), .A2(new_n286), .ZN(new_n637));
  INV_X1    g451(.A(new_n272), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n276), .A2(new_n261), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n295), .B1(new_n641), .B2(new_n317), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n287), .B2(new_n311), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n619), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n414), .A2(new_n415), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT38), .Z(new_n648));
  AND4_X1   g462(.A1(new_n416), .A2(new_n648), .A3(new_n593), .A4(new_n604), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n635), .A2(new_n636), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n421), .ZN(G45));
  INV_X1    g465(.A(new_n629), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n592), .A2(new_n593), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n627), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n315), .A2(new_n575), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n506), .B1(new_n571), .B2(new_n317), .ZN(new_n659));
  AOI211_X1 g473(.A(G469), .B(G902), .C1(new_n568), .C2(new_n570), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n661), .B2(new_n505), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT97), .A4(new_n504), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n571), .A2(new_n317), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G469), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n505), .A3(new_n572), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n658), .A3(new_n505), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT98), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n664), .A2(new_n598), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n315), .A2(new_n671), .A3(new_n351), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  AND3_X1   g488(.A1(new_n664), .A2(new_n609), .A3(new_n670), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n315), .A2(new_n675), .A3(new_n351), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NAND2_X1  g491(.A1(new_n668), .A2(new_n669), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n678), .A2(new_n500), .A3(new_n627), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n315), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  NOR3_X1   g495(.A1(new_n662), .A2(new_n663), .A3(new_n657), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT98), .B1(new_n668), .B2(new_n669), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n290), .A2(new_n291), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n303), .B2(new_n304), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n261), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n303), .A2(new_n686), .A3(new_n304), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n187), .B(KEYINPUT99), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n578), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n596), .A2(new_n593), .A3(new_n604), .A4(new_n607), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n352), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NOR2_X1   g511(.A1(new_n662), .A2(new_n663), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n596), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n692), .A2(new_n578), .A3(new_n619), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n653), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n321), .ZN(G27));
  NAND3_X1  g516(.A1(new_n647), .A2(new_n505), .A3(new_n416), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n533), .B1(new_n532), .B2(new_n534), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n533), .A2(new_n536), .A3(new_n546), .A4(new_n534), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT101), .B(new_n553), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n560), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT101), .B1(new_n549), .B2(new_n553), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n506), .ZN(new_n710));
  NAND2_X1  g524(.A1(G469), .A2(G902), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n572), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n704), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n559), .B1(new_n565), .B2(KEYINPUT101), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n554), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(G469), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(KEYINPUT102), .A3(new_n572), .A4(new_n711), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n653), .B(new_n703), .C1(new_n713), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT104), .B1(new_n311), .B2(new_n287), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n721), .B(KEYINPUT32), .C1(new_n285), .C2(new_n187), .ZN(new_n722));
  INV_X1    g536(.A(new_n279), .ZN(new_n723));
  OAI22_X1  g537(.A1(new_n720), .A2(new_n722), .B1(new_n723), .B2(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n294), .A2(new_n721), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n293), .B1(new_n685), .B2(new_n282), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT103), .B1(new_n726), .B2(KEYINPUT32), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n311), .A2(KEYINPUT104), .A3(new_n287), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n729), .A3(new_n308), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n719), .A2(new_n730), .A3(new_n351), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n352), .B1(new_n310), .B2(new_n314), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n703), .B1(new_n713), .B2(new_n718), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n214), .ZN(G33));
  NOR2_X1   g552(.A1(new_n606), .A2(new_n629), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n315), .A2(new_n351), .A3(new_n739), .A4(new_n734), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n733), .A2(new_n742), .A3(new_n739), .A4(new_n734), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT106), .B(G134), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G36));
  NAND2_X1  g560(.A1(new_n462), .A2(new_n592), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT43), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n613), .A2(new_n748), .A3(new_n620), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n714), .A2(new_n716), .A3(KEYINPUT45), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n752), .B(G469), .C1(KEYINPUT45), .C2(new_n566), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n711), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n572), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n754), .A2(new_n755), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n505), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n595), .B1(new_n414), .B2(new_n415), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT107), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n751), .A2(new_n760), .A3(new_n633), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  INV_X1    g578(.A(new_n761), .ZN(new_n765));
  OR4_X1    g579(.A1(new_n315), .A2(new_n351), .A3(new_n653), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n766), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(G140), .Z(G42));
  OR4_X1    g585(.A1(new_n504), .A2(new_n747), .A3(new_n352), .A4(new_n417), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n661), .B(KEYINPUT108), .Z(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n648), .B(new_n772), .C1(KEYINPUT49), .C2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(new_n645), .C1(KEYINPUT49), .C2(new_n774), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n315), .A2(new_n679), .B1(new_n684), .B2(new_n695), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n672), .A3(new_n676), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n462), .A2(new_n499), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n462), .B2(new_n592), .ZN(new_n781));
  INV_X1    g595(.A(new_n607), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n419), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n575), .A2(new_n613), .A3(new_n351), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n576), .A2(new_n622), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n619), .A2(new_n499), .A3(new_n652), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n603), .A2(new_n461), .A3(new_n605), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n765), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n315), .A2(new_n575), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n700), .A2(new_n653), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n734), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n741), .B2(new_n743), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n732), .A2(new_n736), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n786), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n701), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n713), .A2(new_n718), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n652), .A2(new_n505), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n597), .A2(new_n462), .A3(new_n499), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n644), .A2(new_n620), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n631), .A2(new_n655), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n701), .B1(new_n626), .B2(new_n630), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n655), .A4(new_n801), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT53), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n737), .A2(new_n779), .A3(new_n785), .ZN(new_n809));
  AND4_X1   g623(.A1(KEYINPUT53), .A2(new_n807), .A3(new_n809), .A4(new_n794), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n777), .B(KEYINPUT54), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(new_n807), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n786), .A2(new_n794), .A3(new_n795), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n779), .B(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n737), .A2(new_n812), .A3(new_n785), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n807), .A3(new_n794), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n815), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n811), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT53), .A4(new_n794), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n777), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT111), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n779), .B(KEYINPUT110), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n785), .A2(new_n812), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n794), .A2(new_n795), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n807), .A2(new_n809), .A3(new_n794), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n830), .A2(new_n807), .B1(new_n831), .B2(new_n812), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n824), .A2(new_n777), .B1(new_n832), .B2(new_n820), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n808), .B2(new_n810), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT109), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n730), .A2(new_n351), .ZN(new_n838));
  INV_X1    g652(.A(new_n464), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n748), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n678), .A2(new_n765), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT48), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n464), .A2(new_n645), .A3(new_n351), .A4(new_n841), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n593), .A3(new_n592), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n748), .A2(new_n693), .A3(new_n839), .A4(new_n352), .ZN(new_n846));
  INV_X1    g660(.A(new_n699), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n463), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT115), .Z(new_n850));
  INV_X1    g664(.A(new_n592), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n844), .A2(new_n462), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n841), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n700), .B2(new_n853), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n648), .A2(new_n416), .A3(new_n678), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT113), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n846), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n767), .B(new_n769), .C1(new_n505), .C2(new_n774), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n846), .A2(new_n762), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n862), .B(KEYINPUT51), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n863), .A2(new_n866), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n850), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n826), .A2(new_n837), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n776), .B1(new_n874), .B2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n257), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n832), .A2(new_n317), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n390), .A2(new_n392), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT116), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n398), .B(KEYINPUT55), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n882), .B(new_n883), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n878), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(G51));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n820), .B1(new_n815), .B2(new_n819), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n821), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n711), .B(KEYINPUT57), .Z(new_n892));
  AOI22_X1  g706(.A1(new_n891), .A2(new_n892), .B1(new_n568), .B2(new_n570), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n832), .A2(new_n317), .A3(new_n753), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n888), .B(new_n878), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n821), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n896), .B2(new_n889), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n571), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT117), .B1(new_n898), .B2(new_n877), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n899), .ZN(G54));
  AND2_X1   g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n451), .B1(new_n879), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(KEYINPUT119), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n451), .C1(new_n879), .C2(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n878), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n879), .A2(new_n451), .A3(new_n901), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(G60));
  XNOR2_X1  g724(.A(new_n590), .B(KEYINPUT59), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n891), .A2(new_n588), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n878), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n822), .A2(new_n825), .A3(KEYINPUT111), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n916), .B2(new_n587), .ZN(G63));
  NAND2_X1  g731(.A1(new_n815), .A2(new_n819), .ZN(new_n918));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n617), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n918), .A2(new_n920), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n878), .B(new_n921), .C1(new_n922), .C2(new_n345), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g738(.A(G953), .B1(new_n466), .B2(new_n396), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n786), .B2(G953), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT121), .Z(new_n928));
  OAI21_X1  g742(.A(new_n882), .B1(G898), .B2(new_n257), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(G69));
  XOR2_X1   g744(.A(new_n254), .B(KEYINPUT122), .Z(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n447), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n634), .A2(new_n765), .A3(new_n781), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n733), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n763), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n770), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n650), .A2(new_n655), .A3(new_n805), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n933), .B1(new_n941), .B2(new_n257), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n760), .A2(new_n633), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n838), .A2(new_n593), .A3(new_n604), .A4(new_n596), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n763), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n805), .A2(new_n655), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n946), .A2(new_n770), .A3(new_n737), .A4(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n948), .B2(new_n744), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n257), .A2(G900), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT124), .Z(new_n951));
  OAI21_X1  g765(.A(new_n933), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n943), .A2(new_n955), .A3(new_n953), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n942), .B(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n957), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n960), .B(new_n952), .C1(new_n955), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(G72));
  NOR2_X1   g777(.A1(new_n946), .A2(new_n737), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n770), .A2(new_n947), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n964), .A2(new_n744), .A3(new_n786), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n297), .A2(new_n262), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n877), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n786), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n941), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n262), .A3(new_n297), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n638), .A2(new_n298), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n968), .B(new_n975), .C1(new_n808), .C2(new_n810), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(G57));
endmodule


