//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n202), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G77), .Z(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G244), .Z(new_n222));
  OAI221_X1 g0022(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n226), .B(new_n229), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G226), .B(G232), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n213), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AND2_X1   g0053(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n255));
  OAI21_X1  g0055(.A(G33), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n256), .A2(new_n257), .A3(G68), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT19), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G97), .A2(G107), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n208), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n257), .A2(G33), .A3(G97), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n263), .A2(new_n265), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n230), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT72), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(new_n271), .A3(new_n230), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n260), .A2(new_n267), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g0073(.A(KEYINPUT15), .B(G87), .Z(new_n274));
  NOR2_X1   g0074(.A1(new_n257), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n270), .A2(new_n272), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n274), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n231), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n287), .A2(G244), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n219), .A2(new_n287), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n256), .A2(new_n259), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G116), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n279), .A2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT83), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n294), .A3(G250), .ZN(new_n295));
  AOI21_X1  g0095(.A(G274), .B1(KEYINPUT83), .B2(G250), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n285), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(KEYINPUT69), .A2(G33), .A3(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n231), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n292), .B2(new_n302), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n284), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(G190), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n281), .A2(new_n208), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n273), .A2(new_n310), .A3(new_n277), .ZN(new_n311));
  OAI21_X1  g0111(.A(G200), .B1(new_n292), .B2(new_n302), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT5), .A2(G41), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT5), .A2(G41), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n279), .B(G45), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(new_n301), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G257), .ZN(new_n319));
  OR2_X1    g0119(.A1(KEYINPUT5), .A2(G41), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT5), .A2(G41), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n293), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n301), .A3(G274), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n259), .A2(new_n325), .A3(G250), .A4(G1698), .ZN(new_n326));
  AND2_X1   g0126(.A1(KEYINPUT4), .A2(G244), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n259), .A2(new_n325), .A3(new_n327), .A4(new_n287), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G283), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT4), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n256), .A2(G244), .A3(new_n287), .A4(new_n259), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n319), .B(new_n323), .C1(new_n333), .C2(new_n286), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n306), .ZN(new_n335));
  INV_X1    g0135(.A(new_n286), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n332), .A2(new_n331), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n330), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n338), .A2(new_n304), .A3(new_n319), .A4(new_n323), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G20), .A2(G33), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G77), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n342));
  INV_X1    g0142(.A(G97), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n213), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n264), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n342), .B1(new_n345), .B2(KEYINPUT6), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n259), .A2(new_n325), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(new_n257), .ZN(new_n349));
  OR2_X1    g0149(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n258), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n325), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n349), .B1(new_n353), .B2(KEYINPUT7), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n341), .B(new_n347), .C1(new_n354), .C2(new_n213), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n270), .A2(new_n272), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n276), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n343), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n281), .B2(new_n343), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n335), .B(new_n339), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n355), .B2(new_n356), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n334), .A2(G200), .ZN(new_n363));
  INV_X1    g0163(.A(G190), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n334), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n314), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT8), .B(G58), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n258), .A2(G20), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n369), .B1(G20), .B2(new_n203), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  INV_X1    g0171(.A(new_n340), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n356), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n358), .A2(new_n202), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n356), .B2(new_n358), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n279), .A2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n270), .A2(KEYINPUT73), .A3(new_n272), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n374), .B(new_n375), .C1(new_n380), .C2(new_n202), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n279), .B1(G41), .B2(G45), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n279), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n301), .A2(new_n384), .A3(G274), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT70), .B1(new_n348), .B2(new_n287), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n259), .A2(new_n325), .A3(new_n389), .A4(G1698), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(G223), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n324), .A2(G33), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(G222), .A3(new_n287), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n391), .B(new_n395), .C1(new_n221), .C2(new_n394), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n387), .B1(new_n396), .B2(new_n336), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n301), .A2(G226), .A3(new_n382), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT71), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n381), .B1(new_n403), .B2(G169), .ZN(new_n404));
  AOI21_X1  g0204(.A(G179), .B1(new_n400), .B2(new_n402), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n402), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n401), .B1(new_n397), .B2(new_n398), .ZN(new_n408));
  OAI21_X1  g0208(.A(G190), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT9), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n381), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n381), .A2(KEYINPUT77), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n400), .A2(G200), .A3(new_n402), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n381), .A2(new_n410), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n409), .A2(new_n415), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT10), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n403), .B2(G190), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(new_n416), .A4(new_n415), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n406), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT16), .ZN(new_n425));
  AND2_X1   g0225(.A1(G58), .A2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n426), .B2(new_n201), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n340), .A2(G159), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n427), .A2(KEYINPUT79), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT79), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n254), .A2(new_n255), .A3(G33), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT7), .B(new_n257), .C1(new_n433), .C2(new_n393), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT7), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n394), .B2(G20), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n218), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n425), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(G20), .B1(new_n256), .B2(new_n259), .ZN(new_n439));
  OAI21_X1  g0239(.A(G68), .B1(new_n439), .B2(new_n435), .ZN(new_n440));
  AOI211_X1 g0240(.A(KEYINPUT7), .B(G20), .C1(new_n256), .C2(new_n259), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n431), .B(KEYINPUT16), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n356), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n301), .A2(G232), .A3(new_n382), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n386), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G190), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G226), .A2(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G223), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(G1698), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n256), .A2(new_n259), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n258), .A2(new_n208), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n447), .B1(new_n454), .B2(new_n336), .ZN(new_n455));
  AOI211_X1 g0255(.A(KEYINPUT80), .B(new_n286), .C1(new_n451), .C2(new_n453), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n446), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G200), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n286), .B1(new_n451), .B2(new_n453), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n445), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n368), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n358), .A2(new_n367), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n443), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT17), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n443), .A2(new_n461), .A3(new_n464), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n386), .A2(new_n304), .A3(new_n444), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n455), .B2(new_n456), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n306), .B1(new_n459), .B2(new_n445), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n442), .A2(new_n356), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n434), .A2(new_n436), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G68), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT16), .B1(new_n484), .B2(new_n431), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n464), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT18), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n392), .B1(new_n488), .B2(G33), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n452), .B1(new_n489), .B2(new_n450), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT80), .B1(new_n490), .B2(new_n286), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n459), .A2(new_n447), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n474), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n478), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT81), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n486), .A2(new_n495), .A3(KEYINPUT18), .A4(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n473), .B1(new_n487), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT14), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n301), .A2(G238), .A3(new_n382), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n386), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n212), .A2(new_n287), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n207), .A2(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n259), .A2(new_n503), .A3(new_n325), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n286), .B1(new_n505), .B2(new_n261), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT13), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n506), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT13), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n386), .A4(new_n501), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n500), .B1(new_n511), .B2(G169), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n511), .A2(new_n304), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n500), .A3(G169), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n358), .A2(new_n218), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT12), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n369), .A2(G77), .B1(new_n340), .B2(G50), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n257), .B2(G68), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n356), .A3(KEYINPUT11), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n270), .A2(G68), .A3(new_n272), .A4(new_n378), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n356), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT11), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n519), .A2(new_n522), .A3(new_n523), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n511), .A2(G200), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n507), .A2(new_n510), .A3(G190), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n220), .A2(new_n276), .ZN(new_n533));
  INV_X1    g0333(.A(G77), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n356), .A2(new_n534), .A3(new_n275), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n220), .A2(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n274), .A2(new_n369), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n367), .B(KEYINPUT75), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n372), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n533), .B(new_n535), .C1(new_n539), .C2(new_n356), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n301), .A2(new_n382), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n222), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n388), .A2(G238), .A3(new_n390), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n348), .A2(G107), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n259), .A2(new_n325), .A3(G232), .A4(new_n287), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n543), .A2(new_n544), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n387), .B(new_n542), .C1(new_n549), .C2(new_n336), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n540), .B1(new_n304), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G169), .B2(new_n550), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n528), .A2(new_n532), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n499), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n542), .B1(new_n549), .B2(new_n336), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n458), .B1(new_n555), .B2(new_n386), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n533), .B1(new_n539), .B2(new_n356), .ZN(new_n557));
  INV_X1    g0357(.A(new_n535), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT76), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n550), .A2(G190), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT76), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n540), .C1(new_n550), .C2(new_n458), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n424), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n208), .A2(G20), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n256), .A2(new_n259), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n256), .A2(new_n569), .A3(new_n259), .A4(new_n566), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(KEYINPUT22), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n394), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n369), .A2(G116), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n257), .A2(G107), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n257), .C2(G107), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n579), .A2(new_n580), .B1(new_n578), .B2(new_n577), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n574), .A2(KEYINPUT24), .A3(new_n575), .A4(new_n581), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n356), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n209), .A2(new_n287), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n256), .A2(new_n259), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n336), .B1(new_n318), .B2(G264), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n323), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n458), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G190), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n358), .A2(new_n213), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n282), .B2(G107), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n586), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n214), .A2(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n587), .A2(new_n287), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n256), .A2(new_n259), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(G303), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(new_n394), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n336), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n317), .A2(new_n301), .A3(G270), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n323), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n323), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n282), .A2(G116), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n329), .B(new_n257), .C1(G33), .C2(new_n343), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n248), .A2(G20), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n269), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT20), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n358), .A2(new_n248), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(G169), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n606), .B(G190), .C1(new_n609), .C2(new_n610), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n323), .A2(new_n607), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT84), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n323), .A2(new_n607), .A3(new_n608), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n336), .B2(new_n605), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n623), .B(new_n624), .C1(new_n628), .C2(new_n458), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G179), .A3(new_n619), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n611), .A2(KEYINPUT21), .A3(new_n619), .A4(G169), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n622), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n586), .A2(new_n599), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n594), .A2(G179), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n306), .B2(new_n594), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n366), .A2(new_n565), .A3(new_n600), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n339), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(new_n362), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n314), .A2(new_n639), .A3(KEYINPUT26), .A4(new_n335), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n308), .A2(new_n313), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n361), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n366), .A2(new_n600), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n622), .A2(new_n630), .A3(new_n631), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n633), .B2(new_n635), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n308), .B(new_n644), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n565), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n486), .A2(new_n495), .A3(new_n496), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n497), .ZN(new_n653));
  INV_X1    g0453(.A(new_n552), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n532), .B1(new_n527), .B2(new_n517), .ZN(new_n655));
  INV_X1    g0455(.A(new_n473), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n420), .A2(new_n423), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n406), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n649), .A2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G20), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n279), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n624), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n632), .B2(new_n670), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT87), .Z(new_n673));
  XNOR2_X1  g0473(.A(KEYINPUT88), .B(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n633), .A2(new_n668), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n676), .A2(new_n600), .B1(new_n633), .B2(new_n635), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n633), .A2(new_n635), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n668), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n646), .A2(new_n669), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n679), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n227), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n265), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n233), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n648), .A2(new_n669), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n648), .B2(new_n669), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n636), .A2(new_n366), .A3(new_n600), .A4(new_n669), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n626), .A2(new_n627), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(G179), .A3(new_n303), .A4(new_n606), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n338), .A2(new_n319), .A3(new_n323), .A4(new_n593), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT89), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n334), .A2(new_n304), .ZN(new_n706));
  INV_X1    g0506(.A(new_n303), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n594), .A4(new_n611), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT89), .B(new_n709), .C1(new_n702), .C2(new_n703), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n668), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n700), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n674), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n699), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n694), .B1(new_n719), .B2(G1), .ZN(G364));
  NAND2_X1  g0520(.A1(new_n662), .A2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n690), .A2(G1), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n394), .A2(G355), .A3(new_n227), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n252), .A2(G45), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n489), .A2(new_n688), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G45), .B2(new_n233), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n723), .B1(G116), .B2(new_n227), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  OR3_X1    g0527(.A1(KEYINPUT90), .A2(G13), .A3(G33), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT90), .B1(G13), .B2(G33), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n230), .B1(G20), .B2(new_n306), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n722), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n732), .ZN(new_n736));
  INV_X1    g0536(.A(new_n733), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n257), .A2(new_n364), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n458), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n208), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n304), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n741), .B1(G58), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n304), .A2(new_n458), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n202), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n257), .A2(G190), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n751), .A2(KEYINPUT32), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT32), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n257), .B1(new_n750), .B2(G190), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n753), .B(new_n754), .C1(new_n343), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n749), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n742), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n394), .B1(new_n757), .B2(new_n213), .C1(new_n221), .C2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n748), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n746), .A2(new_n749), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n218), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n740), .A2(new_n604), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n757), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n755), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n394), .B(new_n766), .C1(G294), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n761), .ZN(new_n769));
  INV_X1    g0569(.A(G317), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT33), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(KEYINPUT33), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n747), .B(KEYINPUT91), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G326), .ZN(new_n775));
  INV_X1    g0575(.A(new_n751), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G322), .A2(new_n744), .B1(new_n776), .B2(G329), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n768), .A2(new_n773), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n762), .B1(new_n763), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n735), .B1(new_n672), .B2(new_n736), .C1(new_n737), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n675), .A2(new_n722), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n673), .A2(new_n674), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(G396));
  AOI22_X1  g0585(.A1(G143), .A2(new_n744), .B1(new_n769), .B2(G150), .ZN(new_n786));
  INV_X1    g0586(.A(G137), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n786), .B1(new_n787), .B2(new_n747), .C1(new_n752), .C2(new_n758), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n489), .B1(new_n790), .B2(new_n751), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT94), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n755), .A2(new_n206), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n757), .A2(new_n218), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n789), .B(new_n797), .C1(new_n202), .C2(new_n740), .ZN(new_n798));
  INV_X1    g0598(.A(new_n757), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G87), .A2(new_n799), .B1(new_n776), .B2(G311), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n604), .B2(new_n747), .ZN(new_n801));
  INV_X1    g0601(.A(new_n740), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G107), .B2(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n348), .B1(new_n758), .B2(new_n248), .C1(new_n764), .C2(new_n761), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G97), .B2(new_n767), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n803), .B(new_n805), .C1(new_n806), .C2(new_n743), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n737), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n730), .A2(new_n733), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n722), .B(new_n808), .C1(new_n534), .C2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n552), .A2(new_n668), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n559), .A2(new_n668), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n564), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n552), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n811), .B1(new_n731), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n695), .B(new_n815), .Z(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n717), .ZN(new_n818));
  INV_X1    g0618(.A(new_n722), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(G384));
  INV_X1    g0620(.A(KEYINPUT97), .ZN(new_n821));
  INV_X1    g0621(.A(new_n666), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n486), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n650), .A2(new_n823), .A3(new_n825), .A4(new_n465), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n650), .A2(new_n465), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n499), .A2(new_n824), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n821), .B1(new_n829), .B2(KEYINPUT38), .ZN(new_n830));
  INV_X1    g0630(.A(new_n441), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT7), .B1(new_n489), .B2(G20), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(G68), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT16), .B1(new_n833), .B2(new_n431), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n464), .B1(new_n834), .B2(new_n482), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n822), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n499), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n495), .A3(new_n496), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n839), .A2(new_n465), .A3(new_n836), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n826), .B1(new_n840), .B2(new_n825), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n828), .A2(new_n826), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n823), .B1(new_n653), .B2(new_n473), .ZN(new_n845));
  OAI211_X1 g0645(.A(KEYINPUT97), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n830), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n814), .A2(new_n552), .ZN(new_n848));
  INV_X1    g0648(.A(new_n532), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n527), .B(new_n668), .C1(new_n517), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n527), .A2(new_n668), .ZN(new_n851));
  AOI211_X1 g0651(.A(KEYINPUT14), .B(new_n306), .C1(new_n507), .C2(new_n510), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n512), .A2(new_n852), .A3(new_n514), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n532), .B(new_n851), .C1(new_n853), .C2(new_n529), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n812), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n848), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n716), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g0659(.A1(KEYINPUT100), .A2(KEYINPUT40), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n716), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n847), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT40), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n841), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n838), .B2(new_n841), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n861), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n565), .A2(new_n716), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n674), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT39), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n830), .A2(new_n874), .A3(new_n842), .A4(new_n846), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT98), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT39), .B1(new_n864), .B2(new_n865), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n528), .A2(new_n668), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n648), .A2(new_n669), .A3(new_n815), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n883), .A2(KEYINPUT96), .A3(new_n856), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT96), .B1(new_n883), .B2(new_n856), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n855), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n886), .A2(new_n866), .B1(new_n653), .B2(new_n822), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT99), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n875), .A2(new_n877), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT98), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n880), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n653), .A2(new_n822), .ZN(new_n894));
  INV_X1    g0694(.A(new_n855), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n883), .A2(new_n856), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT96), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n883), .A2(KEYINPUT96), .A3(new_n856), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n894), .B1(new_n900), .B2(new_n867), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n893), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n873), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n565), .B1(new_n696), .B2(new_n698), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n659), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n279), .B2(new_n662), .ZN(new_n908));
  OAI211_X1 g0708(.A(G20), .B(new_n231), .C1(new_n346), .C2(KEYINPUT35), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n248), .B(new_n909), .C1(KEYINPUT35), .C2(new_n346), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT36), .Z(new_n911));
  OAI21_X1  g0711(.A(new_n220), .B1(new_n206), .B2(new_n218), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n912), .A2(new_n233), .B1(G50), .B2(new_n218), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(G1), .A3(new_n661), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(new_n914), .ZN(G367));
  OAI211_X1 g0715(.A(new_n361), .B(new_n365), .C1(new_n362), .C2(new_n669), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n639), .A2(new_n335), .A3(new_n668), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n683), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n680), .A2(new_n685), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n921), .A2(KEYINPUT42), .A3(new_n919), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n361), .B1(new_n678), .B2(new_n916), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n669), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT42), .B1(new_n921), .B2(new_n919), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n311), .A2(new_n669), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n314), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT101), .Z(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n308), .B2(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n920), .A2(new_n932), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT102), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n934), .B2(new_n935), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n689), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n686), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT103), .B1(new_n943), .B2(new_n919), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT103), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n686), .A2(new_n945), .A3(new_n918), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n919), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(KEYINPUT45), .B1(KEYINPUT44), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n946), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n682), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n949), .A2(new_n683), .A3(new_n950), .A4(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n681), .A2(new_n684), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n921), .ZN(new_n958));
  INV_X1    g0758(.A(new_n675), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n719), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n942), .B1(new_n963), .B2(new_n719), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n721), .A2(G1), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n939), .B(new_n940), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n755), .A2(new_n218), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n394), .B1(new_n751), .B2(new_n787), .C1(new_n202), .C2(new_n758), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G58), .C2(new_n802), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n221), .A2(new_n757), .B1(new_n371), .B2(new_n743), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n774), .B2(G143), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n752), .C2(new_n761), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT107), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n757), .A2(new_n343), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G303), .B2(new_n744), .ZN(new_n975));
  INV_X1    g0775(.A(new_n774), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n765), .ZN(new_n977));
  XOR2_X1   g0777(.A(KEYINPUT106), .B(G317), .Z(new_n978));
  AOI211_X1 g0778(.A(new_n489), .B(new_n977), .C1(new_n776), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n802), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n740), .B2(new_n248), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n806), .C2(new_n761), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT105), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n758), .A2(new_n764), .B1(new_n755), .B2(new_n213), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT104), .Z(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n973), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n722), .B1(new_n989), .B2(new_n733), .ZN(new_n990));
  INV_X1    g0790(.A(new_n274), .ZN(new_n991));
  INV_X1    g0791(.A(new_n725), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n734), .B1(new_n227), .B2(new_n991), .C1(new_n243), .C2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n990), .B(new_n993), .C1(new_n736), .C2(new_n930), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n966), .A2(new_n994), .ZN(G387));
  OR2_X1    g0795(.A1(new_n960), .A2(new_n719), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n962), .B1(new_n996), .B2(KEYINPUT109), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n689), .C1(KEYINPUT109), .C2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n960), .A2(new_n965), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT108), .Z(new_n1000));
  INV_X1    g0800(.A(new_n758), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n744), .A2(new_n978), .B1(new_n1001), .B2(G303), .ZN(new_n1002));
  INV_X1    g0802(.A(G322), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n765), .B2(new_n761), .C1(new_n976), .C2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n764), .B2(new_n755), .C1(new_n806), .C2(new_n740), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT49), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n776), .A2(G326), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n489), .B1(G116), .B2(new_n799), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n758), .A2(new_n218), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n761), .A2(new_n367), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n974), .B(new_n1012), .C1(new_n220), .C2(new_n802), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n743), .A2(new_n202), .B1(new_n751), .B2(new_n371), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n747), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(G159), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n767), .A2(new_n274), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n489), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n538), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1020), .A2(G116), .A3(new_n265), .ZN(new_n1021));
  INV_X1    g0821(.A(G45), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(G68), .A2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT50), .B1(new_n538), .B2(G50), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n992), .B1(new_n240), .B2(G45), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n691), .A2(new_n348), .A3(new_n688), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(G107), .B2(new_n227), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1019), .A2(new_n733), .B1(new_n734), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n819), .C1(new_n680), .C2(new_n736), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n998), .A2(new_n1000), .A3(new_n1031), .ZN(G393));
  NAND2_X1  g0832(.A1(new_n955), .A2(new_n956), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n961), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n689), .A3(new_n963), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n955), .A2(new_n965), .A3(new_n956), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n734), .B1(new_n343), .B2(new_n227), .C1(new_n249), .C2(new_n992), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT110), .Z(new_n1038));
  NOR2_X1   g0838(.A1(new_n758), .A2(new_n806), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n761), .A2(new_n604), .B1(new_n751), .B2(new_n1003), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G283), .C2(new_n802), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n747), .A2(new_n770), .B1(new_n743), .B2(new_n765), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT52), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n394), .B1(new_n799), .B2(G107), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n767), .A2(G116), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n538), .A2(new_n758), .B1(new_n202), .B2(new_n761), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT112), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G68), .A2(new_n802), .B1(new_n776), .B2(G143), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT111), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n489), .B1(new_n534), .B2(new_n755), .C1(new_n208), .C2(new_n757), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n747), .A2(new_n371), .B1(new_n743), .B2(new_n752), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n1046), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n722), .B1(new_n1055), .B2(new_n733), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1038), .B(new_n1056), .C1(new_n918), .C2(new_n736), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1035), .A2(new_n1036), .A3(new_n1057), .ZN(G390));
  NAND3_X1  g0858(.A1(new_n857), .A2(new_n716), .A3(G330), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n857), .A2(new_n716), .A3(KEYINPUT113), .A4(G330), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n890), .A2(new_n891), .B1(new_n881), .B2(new_n886), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n896), .A2(new_n855), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n881), .A3(new_n847), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1064), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n878), .A2(new_n879), .B1(new_n900), .B2(new_n880), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n857), .A2(new_n716), .A3(new_n674), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT115), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n716), .A2(G330), .A3(new_n815), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(KEYINPUT114), .A3(new_n895), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n896), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n895), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT114), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1072), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n716), .A2(new_n674), .A3(new_n815), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n895), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1061), .A2(new_n1083), .A3(new_n1062), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n898), .A2(new_n899), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1078), .A2(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n565), .A2(G330), .A3(new_n716), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n905), .A2(new_n1087), .A3(new_n659), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1074), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1088), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(KEYINPUT114), .A2(new_n1071), .B1(new_n1075), .B2(new_n895), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(KEYINPUT115), .B(new_n1090), .C1(new_n1091), .C2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1069), .A2(new_n1073), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT116), .B1(new_n1096), .B2(new_n690), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1065), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1063), .B1(new_n1070), .B2(new_n1067), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1081), .A2(new_n1077), .A3(new_n1076), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT115), .B1(new_n1102), .B2(new_n1090), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1074), .B(new_n1088), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1098), .A2(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n689), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1097), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n965), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n730), .B1(new_n878), .B2(new_n879), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n802), .A2(G150), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1114), .A2(KEYINPUT53), .B1(new_n752), .B2(new_n755), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n348), .B(new_n1115), .C1(KEYINPUT53), .C2(new_n1114), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n776), .A2(G125), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  AOI22_X1  g0918(.A1(new_n769), .A2(G137), .B1(new_n1001), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT117), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n743), .A2(new_n790), .B1(new_n757), .B2(new_n202), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G128), .B2(new_n1015), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G97), .A2(new_n1001), .B1(new_n776), .B2(G294), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n764), .B2(new_n747), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1125), .A2(new_n394), .A3(new_n741), .A4(new_n796), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n743), .A2(new_n248), .B1(new_n755), .B2(new_n534), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT118), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(new_n213), .C2(new_n761), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n737), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n367), .B2(new_n809), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1113), .A2(new_n819), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1111), .A2(new_n1112), .A3(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(KEYINPUT55), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n424), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n424), .A2(new_n1134), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n381), .A2(new_n822), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT56), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OR3_X1    g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n870), .A2(G330), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n862), .A2(KEYINPUT40), .B1(new_n867), .B2(new_n868), .ZN(new_n1145));
  INV_X1    g0945(.A(G330), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n882), .A2(KEYINPUT99), .A3(new_n887), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n893), .B1(new_n892), .B2(new_n901), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n888), .A2(new_n902), .A3(new_n1143), .A4(new_n1147), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n965), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n809), .A2(new_n202), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1015), .A2(G116), .B1(new_n799), .B2(G58), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n764), .B2(new_n751), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G107), .B2(new_n744), .ZN(new_n1157));
  INV_X1    g0957(.A(G41), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n343), .B2(new_n761), .C1(new_n221), .C2(new_n740), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1159), .A2(new_n489), .A3(new_n967), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(new_n1160), .C1(new_n991), .C2(new_n758), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT58), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1158), .B1(new_n488), .B2(new_n258), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n202), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n802), .A2(new_n1118), .B1(new_n1001), .B2(G137), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n744), .A2(G128), .B1(new_n767), .B2(G150), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1015), .A2(G125), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n769), .A2(G132), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G33), .B1(new_n776), .B2(G124), .ZN(new_n1172));
  AOI21_X1  g0972(.A(G41), .B1(new_n799), .B2(G159), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1162), .A2(new_n1164), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n722), .B1(new_n1175), .B2(new_n733), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1154), .B(new_n1176), .C1(new_n1142), .C2(new_n731), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1153), .A2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1152), .B(new_n1151), .C1(new_n1096), .C2(new_n1088), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n689), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1105), .A2(new_n1090), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1178), .B1(new_n1181), .B2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1102), .A2(new_n965), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT120), .Z(new_n1187));
  NOR2_X1   g0987(.A1(new_n747), .A2(new_n806), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n757), .A2(new_n534), .B1(new_n751), .B2(new_n604), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G97), .C2(new_n802), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n348), .B1(new_n761), .B2(new_n248), .C1(new_n764), .C2(new_n743), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n274), .B2(new_n767), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n213), .C2(new_n758), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n747), .A2(new_n790), .B1(new_n758), .B2(new_n371), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n769), .B2(new_n1118), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n489), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G50), .B2(new_n767), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n743), .A2(new_n787), .B1(new_n757), .B2(new_n206), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G159), .B2(new_n802), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n776), .A2(G128), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1197), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n737), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n218), .B2(new_n809), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n819), .B(new_n1203), .C1(new_n855), .C2(new_n731), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1187), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n941), .B(KEYINPUT119), .Z(new_n1207));
  NAND3_X1  g1007(.A1(new_n1109), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(G381));
  AND4_X1   g1009(.A1(new_n1112), .A2(new_n1111), .A3(new_n1178), .A4(new_n1132), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1184), .B2(new_n1181), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(G381), .A2(G393), .A3(G396), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1211), .ZN(G409));
  AOI21_X1  g1016(.A(KEYINPUT122), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT60), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n690), .B1(new_n1108), .B2(new_n1206), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1205), .A2(G384), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G384), .B1(new_n1205), .B2(new_n1220), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n667), .A2(G213), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G375), .B2(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1207), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1179), .B2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1182), .A2(KEYINPUT121), .A3(new_n1183), .A4(new_n1207), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1210), .A2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1228), .A2(new_n1234), .A3(KEYINPUT126), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT126), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1226), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT127), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1228), .A2(new_n1234), .A3(new_n1223), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT123), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT123), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1228), .A2(new_n1234), .A3(new_n1241), .A4(new_n1223), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1225), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n1226), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1238), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1227), .A2(G2897), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1223), .B(new_n1249), .Z(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G390), .A2(new_n966), .A3(new_n994), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(G393), .B(G396), .Z(new_n1258));
  NAND4_X1  g1058(.A1(G390), .A2(new_n966), .A3(KEYINPUT124), .A4(new_n994), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT125), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1257), .A2(new_n1262), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1256), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(new_n1258), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1254), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1252), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1264), .A2(new_n1267), .B1(new_n1270), .B2(new_n1250), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT63), .B(new_n1223), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1243), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1269), .A2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G375), .A2(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1211), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(new_n1224), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1268), .B(new_n1280), .ZN(G402));
endmodule


