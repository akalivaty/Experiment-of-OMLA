//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT69), .A3(KEYINPUT26), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n216), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n210), .B(new_n211), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT66), .B(G190gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT68), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n218), .B1(KEYINPUT28), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n219), .A2(new_n220), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(new_n211), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n211), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n235), .B2(new_n209), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n237), .A3(KEYINPUT25), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g039(.A(G190gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n227), .A2(new_n241), .A3(KEYINPUT64), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n211), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n242), .A2(new_n244), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n240), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n238), .A2(new_n239), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n239), .B1(new_n238), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n226), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G113gat), .B(G120gat), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(new_n256), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n262));
  INV_X1    g061(.A(G134gat), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n263), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n262), .B(new_n264), .C1(KEYINPUT1), .C2(new_n258), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n261), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT25), .B1(new_n237), .B2(new_n248), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT25), .B(new_n233), .C1(new_n235), .C2(new_n209), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n230), .A2(new_n231), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n228), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n238), .A2(new_n250), .A3(new_n239), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n276), .A2(new_n277), .B1(new_n225), .B2(new_n222), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n269), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n208), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n206), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n253), .A2(new_n270), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n269), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n207), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT34), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n283), .A2(new_n284), .A3(new_n287), .A4(new_n207), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n207), .B1(new_n283), .B2(new_n284), .ZN(new_n291));
  INV_X1    g090(.A(new_n281), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n205), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(new_n286), .A3(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n290), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n290), .B2(new_n294), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n202), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n290), .A2(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n295), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n290), .A2(new_n294), .A3(new_n296), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(KEYINPUT36), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT0), .ZN(new_n306));
  XNOR2_X1  g105(.A(G57gat), .B(G85gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G141gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT81), .B(G141gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR3_X1   g114(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n318));
  INV_X1    g117(.A(new_n311), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n310), .A2(G141gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT79), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(G155gat), .B2(G162gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n315), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n321), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n327), .A2(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n317), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n261), .A2(new_n265), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT5), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n331), .A2(new_n332), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n267), .A2(new_n268), .A3(new_n331), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n343), .C1(new_n339), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n317), .B(new_n347), .C1(new_n329), .C2(new_n330), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n332), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n334), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n337), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n349), .B(new_n353), .C1(new_n344), .C2(KEYINPUT4), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n335), .A2(KEYINPUT5), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n309), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  INV_X1    g157(.A(new_n356), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n267), .A2(new_n268), .A3(new_n331), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(KEYINPUT4), .B1(new_n340), .B2(KEYINPUT82), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n350), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n308), .C1(new_n362), .C2(new_n337), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT6), .B(new_n309), .C1(new_n352), .C2(new_n356), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n278), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n226), .B1(new_n272), .B2(new_n275), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n367), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT74), .B(G197gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G204gat), .ZN(new_n374));
  INV_X1    g173(.A(G204gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G197gat), .ZN(new_n377));
  INV_X1    g176(.A(G197gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT74), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G211gat), .A2(G218gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n374), .A2(new_n380), .B1(new_n383), .B2(new_n382), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n391), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n369), .A2(new_n372), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n367), .B1(new_n278), .B2(KEYINPUT29), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n250), .A2(new_n238), .B1(new_n222), .B2(new_n225), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n367), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n368), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G8gat), .B(G36gat), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT78), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n368), .B1(new_n253), .B2(new_n371), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n401), .A2(new_n400), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n372), .B1(new_n253), .B2(new_n367), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n403), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT30), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n409), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n411), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n366), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n426), .B(KEYINPUT83), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT86), .B(G22gat), .ZN(new_n429));
  INV_X1    g228(.A(G228gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n348), .A2(new_n371), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n395), .A2(new_n392), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n385), .A2(new_n387), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n371), .B1(new_n389), .B2(new_n386), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n347), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n331), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n432), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n432), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n347), .B1(new_n393), .B2(KEYINPUT29), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n331), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n433), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n404), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n433), .A2(new_n445), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n429), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n439), .A2(new_n440), .ZN(new_n451));
  AOI211_X1 g250(.A(KEYINPUT84), .B(new_n432), .C1(new_n434), .C2(new_n438), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n449), .B(new_n429), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n428), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G22gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n453), .A3(new_n426), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n423), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n458), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n354), .A2(new_n335), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT39), .C1(new_n335), .C2(new_n333), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n354), .A2(new_n463), .A3(new_n335), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(new_n308), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n464), .B2(new_n308), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n411), .A2(new_n419), .A3(new_n421), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT40), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n357), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n460), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n415), .B2(new_n404), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT88), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT38), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n409), .B1(new_n420), .B2(KEYINPUT37), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n417), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n410), .B1(new_n405), .B2(new_n475), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n420), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n485), .A2(new_n366), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n304), .B(new_n459), .C1(new_n474), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n297), .A2(new_n298), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n460), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n494), .B2(new_n423), .ZN(new_n495));
  INV_X1    g294(.A(new_n423), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n460), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(G71gat), .A2(G78gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n501));
  NAND2_X1  g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT100), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(G57gat), .A2(G64gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n503), .A2(new_n506), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT99), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  INV_X1    g313(.A(G57gat), .ZN(new_n515));
  INV_X1    g314(.A(G64gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT99), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n514), .A2(new_n519), .A3(new_n508), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n500), .A2(new_n521), .A3(new_n502), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT98), .B1(new_n504), .B2(new_n505), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n512), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G127gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(G1gat), .B2(new_n532), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G8gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(new_n526), .B2(new_n525), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n531), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n322), .ZN(new_n541));
  XOR2_X1   g340(.A(G183gat), .B(G211gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n539), .B(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(KEYINPUT41), .ZN(new_n546));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT92), .B(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G36gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT92), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G36gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT93), .A3(G29gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G43gat), .A2(G50gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT15), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(G43gat), .ZN(new_n565));
  INV_X1    g364(.A(G50gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n561), .ZN(new_n569));
  NOR2_X1   g368(.A1(G29gat), .A2(G36gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n570), .A2(new_n574), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n564), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n578));
  NOR2_X1   g377(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n578), .A2(new_n579), .B1(G29gat), .B2(G36gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n574), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n580), .A2(new_n581), .B1(new_n558), .B2(G29gat), .ZN(new_n582));
  OAI22_X1  g381(.A1(new_n560), .A2(new_n577), .B1(new_n582), .B2(new_n564), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT94), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  OAI221_X1 g384(.A(new_n585), .B1(new_n582), .B2(new_n564), .C1(new_n560), .C2(new_n577), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n584), .A2(new_n586), .A3(new_n590), .A4(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n593), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n596), .A2(new_n600), .A3(new_n603), .A4(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n609));
  OR3_X1    g408(.A1(new_n583), .A2(new_n609), .A3(new_n587), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n583), .B2(new_n587), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n584), .A2(new_n586), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n614), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n545), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n613), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n549), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n548), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n525), .A2(new_n607), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n514), .A2(new_n519), .A3(new_n508), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n523), .A3(new_n522), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n628), .A2(new_n512), .A3(new_n606), .A4(new_n605), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n512), .A4(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(KEYINPUT102), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n544), .A2(new_n624), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT90), .B(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT11), .B(G169gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n536), .B1(new_n610), .B2(new_n611), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n592), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n614), .A2(new_n536), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT18), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n656), .A2(new_n657), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n657), .B(KEYINPUT13), .Z(new_n664));
  NOR2_X1   g463(.A1(new_n614), .A2(new_n536), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n658), .B1(new_n592), .B2(new_n655), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n662), .B1(new_n668), .B2(new_n657), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n654), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n661), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n672), .A2(new_n663), .A3(new_n666), .A4(new_n653), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n647), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n499), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n366), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g479(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n471), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT104), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(G8gat), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n688));
  OAI22_X1  g487(.A1(new_n684), .A2(new_n687), .B1(new_n682), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(new_n677), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n690), .B2(new_n304), .ZN(new_n691));
  INV_X1    g490(.A(new_n493), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n693), .ZN(G1326gat));
  INV_X1    g493(.A(new_n460), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT105), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n624), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n499), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n646), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n675), .A2(new_n544), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n552), .A3(new_n678), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n701), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n712));
  NAND3_X1  g511(.A1(new_n499), .A2(new_n700), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n704), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT107), .B1(new_n715), .B2(new_n366), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n366), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n707), .B1(new_n717), .B2(new_n718), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n422), .A2(new_n558), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n551), .B1(new_n714), .B2(new_n471), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n722), .B(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n724), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(new_n304), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G43gat), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n701), .A2(new_n692), .A3(new_n704), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n715), .A2(new_n732), .B1(G43gat), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g534(.A(new_n566), .B1(new_n714), .B2(new_n695), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n695), .A2(new_n566), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT109), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n705), .A2(new_n739), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n737), .B1(new_n736), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1331gat));
  INV_X1    g542(.A(new_n544), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n744), .A2(new_n674), .A3(new_n700), .A4(new_n646), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n499), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n678), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n471), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT49), .B(G64gat), .Z(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(G1333gat));
  NAND2_X1  g551(.A1(new_n746), .A2(new_n731), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n692), .A2(G71gat), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n753), .A2(G71gat), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n746), .A2(new_n695), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n544), .A2(new_n674), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n499), .A2(new_n700), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n499), .A2(KEYINPUT51), .A3(new_n700), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n764), .A2(new_n598), .A3(new_n678), .A4(new_n702), .ZN(new_n765));
  INV_X1    g564(.A(new_n759), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n646), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n711), .B2(new_n713), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n678), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n765), .B1(new_n770), .B2(new_n598), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT110), .B(new_n765), .C1(new_n770), .C2(new_n598), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n499), .A2(new_n700), .A3(new_n712), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n709), .B1(new_n499), .B2(new_n700), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n471), .B(new_n767), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n422), .A2(G92gat), .A3(new_n646), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n776), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n779), .A2(G92gat), .B1(new_n764), .B2(new_n781), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n776), .B1(new_n785), .B2(new_n783), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  INV_X1    g588(.A(G99gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n769), .A2(new_n731), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n764), .A2(new_n790), .A3(new_n493), .A4(new_n702), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n695), .A2(G106gat), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n769), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n460), .A2(new_n646), .ZN(new_n800));
  AOI21_X1  g599(.A(G106gat), .B1(new_n764), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n797), .B(KEYINPUT53), .C1(new_n799), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n769), .B2(new_n798), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n764), .A2(new_n800), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(G106gat), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n802), .A2(new_n807), .ZN(G1339gat));
  NOR2_X1   g607(.A1(new_n675), .A2(G113gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n647), .A2(new_n674), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n658), .A2(new_n665), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n657), .A2(new_n668), .B1(new_n811), .B2(new_n664), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n652), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n673), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT115), .A4(new_n636), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n634), .A3(KEYINPUT54), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n636), .B1(new_n630), .B2(new_n631), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n821));
  AOI21_X1  g620(.A(new_n642), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n634), .A2(new_n637), .A3(new_n642), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT55), .B1(new_n819), .B2(new_n822), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n700), .A2(new_n814), .A3(new_n829), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n702), .A2(new_n814), .B1(new_n829), .B2(new_n674), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n700), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n810), .B1(new_n832), .B2(new_n744), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n366), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n494), .A2(new_n471), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n809), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n836), .B2(new_n675), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1340gat));
  AND2_X1   g641(.A1(new_n834), .A2(new_n835), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g644(.A(G120gat), .B(new_n646), .C1(new_n845), .C2(new_n837), .ZN(new_n846));
  INV_X1    g645(.A(G120gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n843), .B2(new_n702), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n847), .B(new_n702), .C1(new_n838), .C2(new_n839), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  INV_X1    g650(.A(new_n848), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n843), .A2(new_n544), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n530), .A2(KEYINPUT120), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(G1342gat));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n700), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(G134gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n843), .A2(KEYINPUT121), .A3(new_n263), .A4(new_n700), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n859), .A2(G134gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n731), .A2(new_n460), .A3(new_n471), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n834), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(G141gat), .A3(new_n675), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n829), .A2(new_n674), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n673), .A2(new_n813), .A3(new_n702), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n700), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n700), .A2(new_n814), .A3(new_n829), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n744), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n810), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n460), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n879), .B(new_n880), .C1(new_n833), .C2(new_n460), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n823), .A2(new_n825), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n828), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n674), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n673), .A2(new_n813), .A3(new_n702), .A4(KEYINPUT123), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n624), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n544), .B1(new_n889), .B2(new_n830), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n695), .C1(new_n890), .C2(new_n810), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n878), .A2(new_n881), .A3(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n731), .A2(new_n366), .A3(new_n471), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n674), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n870), .B1(new_n894), .B2(new_n312), .ZN(new_n895));
  XNOR2_X1  g694(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n895), .B(new_n897), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n702), .A3(new_n893), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n310), .A2(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT57), .B1(new_n833), .B2(new_n460), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n460), .A2(KEYINPUT57), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n827), .A2(new_n828), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n906), .B2(new_n624), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n700), .A2(new_n829), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n909), .A3(new_n814), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n544), .B1(new_n889), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n911), .B2(new_n810), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n902), .A2(new_n702), .A3(new_n912), .A4(new_n893), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G148gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT59), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n901), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n869), .A2(G148gat), .A3(new_n646), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n899), .A2(new_n900), .B1(new_n914), .B2(KEYINPUT59), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(new_n921), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1345gat));
  INV_X1    g722(.A(new_n869), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n322), .A3(new_n544), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n892), .A2(new_n893), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n544), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(new_n322), .ZN(G1346gat));
  AOI21_X1  g727(.A(G162gat), .B1(new_n924), .B2(new_n700), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n624), .A2(new_n323), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n833), .A2(new_n678), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n494), .A2(new_n422), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n675), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(new_n213), .ZN(G1348gat));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n646), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(new_n214), .ZN(G1349gat));
  NAND3_X1  g737(.A1(new_n932), .A2(new_n544), .A3(new_n933), .ZN(new_n939));
  MUX2_X1   g738(.A(new_n220), .B(G183gat), .S(new_n939), .Z(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g740(.A1(new_n934), .A2(new_n624), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n241), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n219), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1351gat));
  AND2_X1   g746(.A1(new_n902), .A2(new_n912), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n731), .A2(new_n678), .A3(new_n422), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(new_n378), .A3(new_n675), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n932), .A2(new_n695), .A3(new_n471), .A4(new_n304), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n674), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(new_n378), .ZN(G1352gat));
  NOR3_X1   g755(.A1(new_n952), .A2(G204gat), .A3(new_n646), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n948), .A2(new_n702), .A3(new_n949), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n375), .B2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n948), .A2(new_n544), .A3(new_n949), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n953), .A2(new_n954), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n744), .A2(G211gat), .ZN(new_n965));
  OAI22_X1  g764(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n950), .B2(new_n624), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n624), .A2(G218gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n964), .B2(new_n968), .ZN(G1355gat));
endmodule


