//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT68), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT70), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n465), .A3(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(KEYINPUT71), .A3(G136), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n472), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n464), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n479), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n482), .A2(new_n486), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n483), .A2(new_n479), .A3(new_n464), .A4(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n479), .A2(G102), .A3(G2104), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n479), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n475), .B2(G126), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n495), .B(new_n499), .C1(new_n502), .C2(new_n479), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .A3(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  INV_X1    g097(.A(new_n520), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G62), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  NOR2_X1   g101(.A1(new_n516), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n521), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(G52), .A2(new_n527), .B1(new_n521), .B2(G90), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n520), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n527), .A2(G43), .B1(G651), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n521), .A2(G81), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n512), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n521), .A2(G91), .B1(G651), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n527), .A2(KEYINPUT9), .A3(G53), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n527), .A2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n521), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n520), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n510), .A2(G48), .A3(G543), .A4(new_n511), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n523), .A2(new_n510), .A3(G86), .A4(new_n511), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n521), .A2(G85), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n527), .A2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n506), .C2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT74), .Z(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n520), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT75), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G299), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n595), .B2(G168), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(new_n595), .B2(G168), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  OR2_X1    g175(.A1(new_n549), .A2(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n591), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n485), .A2(G123), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n481), .A2(G135), .ZN(new_n606));
  NOR2_X1   g181(.A1(G99), .A2(G2105), .ZN(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(new_n479), .B2(G111), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(G2096), .Z(new_n610));
  NAND3_X1  g185(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT76), .Z(G156));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2435), .ZN(new_n618));
  XOR2_X1   g193(.A(G2427), .B(G2438), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT14), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT77), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT79), .Z(new_n631));
  INV_X1    g206(.A(G14), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n627), .B2(new_n629), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(G401));
  XOR2_X1   g210(.A(G2067), .B(G2678), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n639), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT17), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n640), .A2(new_n644), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n648), .B1(KEYINPUT81), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(KEYINPUT81), .B2(new_n650), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n647), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n655), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n665), .C1(new_n663), .C2(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(G229));
  NOR2_X1   g248(.A1(G5), .A2(G16), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(G301), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1961), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G33), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT25), .Z(new_n685));
  INV_X1    g260(.A(G139), .ZN(new_n686));
  INV_X1    g261(.A(G127), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n467), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G115), .B2(G2104), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n685), .B1(new_n686), .B2(new_n480), .C1(new_n689), .C2(new_n479), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n683), .B1(new_n690), .B2(G29), .ZN(new_n691));
  INV_X1    g266(.A(G2072), .ZN(new_n692));
  INV_X1    g267(.A(G2084), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n682), .B1(new_n694), .B2(G34), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(G34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n477), .B2(new_n682), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n691), .A2(new_n692), .B1(new_n693), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT30), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G28), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G28), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n704), .A3(new_n682), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(G164), .A2(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G27), .B2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G2078), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n708), .A2(new_n709), .B1(new_n691), .B2(new_n692), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n681), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n682), .A2(G35), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n682), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G2090), .ZN(new_n716));
  NAND2_X1  g291(.A1(G299), .A2(G16), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n676), .A2(KEYINPUT23), .A3(G20), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n719));
  INV_X1    g294(.A(G20), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1956), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n712), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n715), .A2(G2090), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n676), .A2(G4), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n592), .B2(new_n676), .ZN(new_n731));
  INV_X1    g306(.A(G1348), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n682), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n481), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n485), .A2(G128), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n479), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(new_n682), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n727), .A2(new_n729), .A3(new_n733), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n676), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n549), .B2(new_n676), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G286), .A2(new_n676), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n753), .B1(new_n752), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G1966), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT92), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n677), .A2(new_n678), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G1966), .B2(new_n756), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n747), .A2(new_n751), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n481), .A2(G131), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n485), .A2(G119), .ZN(new_n763));
  NOR2_X1   g338(.A1(G95), .A2(G2105), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(new_n479), .B2(G107), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G25), .B(new_n766), .S(G29), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT35), .B(G1991), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n676), .A2(G24), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G290), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1986), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n767), .A2(new_n768), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT85), .B1(new_n777), .B2(G16), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n777), .A2(KEYINPUT85), .A3(G16), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n778), .B(new_n779), .C1(G166), .C2(new_n676), .ZN(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G23), .B(G288), .S(G16), .Z(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(new_n791), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n776), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(KEYINPUT86), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT87), .ZN(new_n796));
  AOI21_X1  g371(.A(KEYINPUT86), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n481), .A2(G141), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n485), .A2(G129), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n479), .A2(G105), .A3(G2104), .ZN(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT26), .Z(new_n805));
  NAND4_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G29), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G29), .B2(G32), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n709), .B2(new_n708), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n761), .A2(new_n799), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n700), .A2(new_n693), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n609), .A2(new_n682), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n809), .A2(new_n810), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(G311));
  AND4_X1   g394(.A1(new_n799), .A2(new_n761), .A3(new_n800), .A4(new_n813), .ZN(new_n820));
  INV_X1    g395(.A(new_n815), .ZN(new_n821));
  INV_X1    g396(.A(new_n816), .ZN(new_n822));
  INV_X1    g397(.A(new_n818), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(G150));
  NAND2_X1  g399(.A1(new_n521), .A2(G93), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT95), .B(G55), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n825), .B1(new_n506), .B2(new_n826), .C1(new_n557), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n549), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n599), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT96), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n609), .B(new_n806), .ZN(new_n839));
  INV_X1    g414(.A(G142), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n479), .A2(G118), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n480), .A2(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G130), .B2(new_n485), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n839), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n741), .B(new_n503), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n612), .B(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n846), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n766), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n492), .B(G160), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT100), .B(G37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g433(.A1(new_n828), .A2(new_n595), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n602), .B(new_n829), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n591), .B(G299), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n862), .B(KEYINPUT41), .Z(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n861), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n864), .B(new_n860), .S(new_n866), .Z(new_n867));
  XOR2_X1   g442(.A(G166), .B(G288), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(G305), .ZN(new_n869));
  XOR2_X1   g444(.A(G290), .B(KEYINPUT102), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT42), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n873), .B2(new_n595), .ZN(G295));
  OAI21_X1  g449(.A(new_n859), .B1(new_n873), .B2(new_n595), .ZN(G331));
  XNOR2_X1  g450(.A(new_n829), .B(G286), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G171), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n877), .A2(new_n865), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n863), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n878), .A2(new_n879), .A3(new_n871), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n856), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n880), .A2(new_n884), .A3(new_n885), .A4(new_n881), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(KEYINPUT44), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n884), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n880), .A2(KEYINPUT43), .A3(new_n885), .A4(new_n881), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(G397));
  INV_X1    g467(.A(KEYINPUT126), .ZN(new_n893));
  INV_X1    g468(.A(G1384), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n483), .A2(G126), .A3(new_n464), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n479), .B1(new_n895), .B2(new_n500), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n499), .A2(new_n495), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(G40), .B(new_n470), .C1(new_n476), .C2(G2105), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n741), .B(G2067), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT104), .ZN(new_n905));
  INV_X1    g480(.A(G1996), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n806), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n766), .B(new_n768), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT105), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G290), .B(new_n772), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G8), .ZN(new_n914));
  NOR2_X1   g489(.A1(G166), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT55), .Z(new_n916));
  INV_X1    g491(.A(KEYINPUT50), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n503), .A2(new_n917), .A3(new_n894), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n503), .B2(new_n894), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n901), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n898), .A2(KEYINPUT50), .ZN(new_n923));
  INV_X1    g498(.A(new_n901), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT108), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n919), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(KEYINPUT106), .B(G2090), .Z(new_n927));
  NAND3_X1  g502(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n894), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n900), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n926), .A2(new_n927), .B1(new_n781), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n916), .B1(new_n930), .B2(new_n914), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n781), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n901), .B1(new_n898), .B2(KEYINPUT50), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n918), .A3(new_n927), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n915), .B(KEYINPUT55), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n937), .A2(new_n938), .A3(G8), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n895), .A2(new_n500), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G2105), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n499), .A2(new_n495), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n914), .B1(new_n944), .B2(new_n924), .ZN(new_n945));
  NAND2_X1  g520(.A1(G305), .A2(G1981), .ZN(new_n946));
  INV_X1    g521(.A(G1981), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n574), .A2(new_n576), .A3(new_n947), .A4(new_n575), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(KEYINPUT49), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n945), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n567), .A2(new_n568), .A3(G1976), .A4(new_n569), .ZN(new_n954));
  INV_X1    g529(.A(G1976), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT52), .B1(G288), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n945), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n954), .B(G8), .C1(new_n898), .C2(new_n901), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT52), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT109), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n957), .A3(new_n959), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n931), .A2(new_n940), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n923), .A2(new_n924), .A3(new_n918), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n933), .A2(KEYINPUT111), .A3(new_n918), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n678), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n900), .A2(new_n924), .A3(new_n928), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(KEYINPUT53), .A3(new_n709), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n929), .B2(G2078), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G171), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT119), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT119), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(G171), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(G286), .A2(G8), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT116), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n971), .A2(G1966), .B1(G2084), .B2(new_n966), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(G8), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n985), .A2(KEYINPUT117), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n982), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT62), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n984), .B(G8), .C1(KEYINPUT117), .C2(new_n985), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n986), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n965), .A2(new_n980), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT123), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n986), .A2(new_n989), .A3(new_n991), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT123), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n965), .A2(new_n980), .A3(new_n997), .A4(new_n992), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n940), .ZN(new_n1000));
  INV_X1    g575(.A(new_n960), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n953), .A2(new_n955), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n948), .B1(new_n1002), .B2(G288), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1000), .A2(new_n1001), .B1(new_n1003), .B2(new_n945), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT63), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n932), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT107), .B1(new_n932), .B2(new_n934), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n914), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1008), .B2(new_n938), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1005), .B1(new_n1009), .B2(KEYINPUT110), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n987), .A2(G286), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n1001), .C1(new_n1008), .C2(new_n938), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1010), .A2(new_n940), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n965), .A2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1005), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n999), .A2(new_n1004), .A3(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT56), .B(G2072), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n971), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n926), .B2(G1956), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G299), .B(KEYINPUT57), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(new_n1020), .C1(new_n926), .C2(G1956), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n591), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n968), .A2(new_n732), .A3(new_n969), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  INV_X1    g604(.A(G2067), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n944), .A2(new_n924), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1023), .B1(new_n1027), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT60), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1041), .A3(new_n592), .ZN(new_n1042));
  OAI211_X1 g617(.A(KEYINPUT60), .B(new_n591), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n898), .B2(new_n901), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT113), .B(new_n1045), .C1(new_n898), .C2(new_n901), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n1049), .C1(new_n929), .C2(G1996), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n549), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT59), .B1(new_n1051), .B2(KEYINPUT114), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(KEYINPUT114), .A3(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT61), .A3(new_n1025), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1035), .B1(new_n1044), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g638(.A(new_n979), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n978), .B1(new_n975), .B2(G171), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n971), .A2(new_n1066), .A3(KEYINPUT53), .A4(new_n709), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n971), .A2(KEYINPUT120), .A3(G2078), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n970), .A2(new_n1067), .A3(new_n974), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n974), .A2(G301), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1064), .A2(new_n1065), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT121), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1073), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1075), .B(new_n1076), .C1(new_n980), .C2(new_n1071), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n995), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1069), .A2(G171), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT122), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n975), .A2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1069), .A2(new_n1082), .A3(G171), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(KEYINPUT54), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n965), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1035), .C1(new_n1044), .C2(new_n1061), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1063), .A2(new_n1078), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n913), .B1(new_n1018), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n903), .B1(new_n905), .B2(new_n807), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT46), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(KEYINPUT124), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n902), .A2(new_n906), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(KEYINPUT124), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT47), .Z(new_n1098));
  NOR3_X1   g673(.A1(new_n903), .A2(G1986), .A3(G290), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1100));
  XNOR2_X1  g675(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n911), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n902), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n908), .A2(new_n768), .A3(new_n766), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n742), .A2(new_n1030), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n903), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1098), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n893), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n999), .A2(new_n1017), .A3(new_n1004), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1088), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1059), .A2(KEYINPUT61), .A3(new_n1025), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT61), .B1(new_n1059), .B2(new_n1025), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(new_n1042), .A3(new_n1043), .A4(new_n1056), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1087), .B1(new_n1115), .B2(new_n1035), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n995), .B(new_n1085), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1110), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(KEYINPUT126), .B(new_n1107), .C1(new_n1119), .C2(new_n913), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1109), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g696(.A(G227), .ZN(new_n1123));
  NAND3_X1  g697(.A1(new_n634), .A2(G319), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g698(.A1(new_n1124), .A2(KEYINPUT127), .ZN(new_n1125));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n1126));
  NAND4_X1  g700(.A1(new_n634), .A2(new_n1126), .A3(G319), .A4(new_n1123), .ZN(new_n1127));
  AOI21_X1  g701(.A(G229), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g702(.A1(new_n1128), .A2(new_n857), .A3(new_n888), .A4(new_n889), .ZN(G225));
  INV_X1    g703(.A(G225), .ZN(G308));
endmodule


