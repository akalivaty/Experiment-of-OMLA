//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n655, new_n658, new_n660, new_n661,
    new_n662, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT65), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n461), .A2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G125), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n469), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n466), .A2(KEYINPUT66), .B1(G113), .B2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(new_n476), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n462), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G101), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n489), .B2(G101), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT3), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n461), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n492), .B1(G137), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G160));
  NAND2_X1  g073(.A1(new_n495), .A2(G136), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n480), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G124), .ZN(new_n501));
  OR2_X1    g076(.A1(G100), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n499), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n506), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(G2105), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n493), .A2(new_n461), .A3(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n474), .A2(new_n507), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n480), .A2(G114), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT70), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(new_n511), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n493), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n507), .B1(new_n464), .B2(new_n465), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G164));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT72), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n529), .B1(new_n534), .B2(KEYINPUT6), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n536), .A2(KEYINPUT5), .A3(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(G543), .B1(new_n536), .B2(KEYINPUT5), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G88), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G50), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n542), .B1(new_n545), .B2(KEYINPUT73), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n536), .A2(KEYINPUT5), .A3(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(G62), .ZN(new_n549));
  NAND2_X1  g124(.A1(G75), .A2(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n534), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n541), .A2(new_n544), .A3(new_n552), .ZN(G303));
  INV_X1    g128(.A(G303), .ZN(G166));
  OAI21_X1  g129(.A(KEYINPUT76), .B1(new_n535), .B2(new_n542), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n531), .B2(new_n533), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(G543), .C1(new_n558), .C2(new_n529), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G51), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n540), .A2(G89), .ZN(new_n562));
  NAND3_X1  g137(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT7), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n565), .B1(new_n537), .B2(new_n538), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n547), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(G63), .A3(G651), .A4(new_n567), .ZN(new_n568));
  AND4_X1   g143(.A1(new_n561), .A2(new_n562), .A3(new_n564), .A4(new_n568), .ZN(G168));
  NAND2_X1  g144(.A1(G77), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  INV_X1    g146(.A(G64), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(new_n534), .B1(G90), .B2(new_n540), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n560), .A2(G52), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G301));
  INV_X1    g151(.A(G301), .ZN(G171));
  NAND2_X1  g152(.A1(G68), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G56), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(new_n534), .B1(G81), .B2(new_n540), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n560), .A2(G43), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G860), .ZN(G153));
  NAND4_X1  g160(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g161(.A1(G1), .A2(G3), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT8), .ZN(new_n588));
  NAND4_X1  g163(.A1(G319), .A2(G483), .A3(G661), .A4(new_n588), .ZN(G188));
  INV_X1    g164(.A(G53), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n543), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n543), .B(new_n591), .C1(KEYINPUT77), .C2(KEYINPUT9), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n548), .A2(G65), .ZN(new_n596));
  AND2_X1   g171(.A1(G78), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n540), .A2(G91), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n598), .A4(new_n599), .ZN(G299));
  INV_X1    g175(.A(G168), .ZN(G286));
  INV_X1    g176(.A(G74), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n547), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT75), .B1(new_n546), .B2(new_n547), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  OAI211_X1 g181(.A(G87), .B(new_n548), .C1(new_n558), .C2(new_n529), .ZN(new_n607));
  OAI211_X1 g182(.A(G49), .B(G543), .C1(new_n558), .C2(new_n529), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G288));
  NAND2_X1  g184(.A1(G48), .A2(G543), .ZN(new_n610));
  OR3_X1    g185(.A1(new_n535), .A2(KEYINPUT78), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT78), .B1(new_n535), .B2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(G73), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G61), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n539), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n540), .A2(G86), .B1(new_n616), .B2(new_n534), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G305));
  XNOR2_X1  g193(.A(KEYINPUT72), .B(G651), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n566), .A2(G60), .A3(new_n567), .ZN(new_n620));
  AND2_X1   g195(.A1(G72), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT79), .ZN(new_n624));
  INV_X1    g199(.A(G47), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n555), .B2(new_n559), .ZN(new_n626));
  INV_X1    g201(.A(new_n529), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n619), .B2(new_n557), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n628), .A2(G85), .A3(new_n548), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(KEYINPUT80), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n559), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n556), .B1(new_n628), .B2(G543), .ZN(new_n633));
  OAI21_X1  g208(.A(G47), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT80), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(new_n635), .A3(new_n629), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n624), .A2(new_n631), .A3(new_n636), .ZN(G290));
  INV_X1    g212(.A(G868), .ZN(new_n638));
  NOR2_X1   g213(.A1(G301), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n628), .A2(new_n548), .ZN(new_n642));
  INV_X1    g217(.A(G92), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(G79), .A2(G543), .ZN(new_n645));
  INV_X1    g220(.A(G66), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n539), .B2(new_n646), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n640), .A2(new_n644), .B1(G651), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n560), .A2(G54), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n639), .B1(new_n652), .B2(new_n638), .ZN(G284));
  AOI21_X1  g228(.A(new_n639), .B1(new_n652), .B2(new_n638), .ZN(G321));
  NAND2_X1  g229(.A1(G299), .A2(new_n638), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(G168), .B2(new_n638), .ZN(G297));
  OAI21_X1  g231(.A(new_n655), .B1(G168), .B2(new_n638), .ZN(G280));
  INV_X1    g232(.A(G559), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n658), .B2(G860), .ZN(G148));
  NAND2_X1  g234(.A1(new_n583), .A2(new_n638), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n650), .B(KEYINPUT81), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n661), .A2(G559), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n662), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g238(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g239(.A1(new_n474), .A2(new_n489), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT13), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n495), .A2(G135), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n500), .A2(G123), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n672), .A2(new_n480), .A3(G111), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n480), .B2(G111), .ZN(new_n674));
  OR2_X1    g249(.A1(G99), .A2(G2105), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(G2104), .A3(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n670), .B(new_n671), .C1(new_n673), .C2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT84), .B(G2096), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n669), .A2(new_n679), .ZN(G156));
  XNOR2_X1  g255(.A(G2427), .B(G2438), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2430), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT15), .B(G2435), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(KEYINPUT14), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT86), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1341), .B(G1348), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2451), .B(G2454), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2443), .B(G2446), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n695), .A2(new_n696), .A3(G14), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G401));
  XOR2_X1   g273(.A(G2084), .B(G2090), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G2072), .A2(G2078), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n442), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G2067), .B(G2678), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT18), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n702), .A2(KEYINPUT87), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(KEYINPUT87), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n708), .A3(new_n704), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n702), .B(KEYINPUT17), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n709), .B(new_n700), .C1(new_n710), .C2(new_n704), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n704), .A3(new_n699), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n706), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(G2096), .B(G2100), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(G227));
  XOR2_X1   g290(.A(G1971), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT19), .ZN(new_n717));
  XOR2_X1   g292(.A(G1956), .B(G2474), .Z(new_n718));
  XOR2_X1   g293(.A(G1961), .B(G1966), .Z(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT20), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n718), .A2(new_n719), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n717), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n717), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT88), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(G1991), .B(G1996), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(G1981), .B(G1986), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(G229));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT97), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G139), .B2(new_n495), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(new_n480), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2072), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT30), .B(G28), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n677), .A2(new_n734), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n745), .B1(G29), .B2(new_n746), .C1(new_n747), .C2(KEYINPUT102), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(KEYINPUT102), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G1966), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NOR2_X1   g327(.A1(G168), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(G21), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n751), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT101), .Z(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n755), .A2(new_n757), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n489), .A2(G105), .ZN(new_n763));
  INV_X1    g338(.A(new_n495), .ZN(new_n764));
  INV_X1    g339(.A(G141), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n500), .A2(G129), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n734), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n734), .B2(G32), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT27), .ZN(new_n777));
  INV_X1    g352(.A(G1996), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n762), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT93), .Z(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n652), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n734), .B1(KEYINPUT24), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(KEYINPUT24), .B2(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n497), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n734), .A2(G26), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT28), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n500), .A2(G128), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n480), .A2(G116), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n495), .A2(G140), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n794), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n752), .A2(G5), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G171), .B2(new_n752), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n752), .A2(G19), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n583), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT95), .B(G1341), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n804), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n734), .A2(G35), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G162), .B2(new_n734), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT29), .Z(new_n817));
  INV_X1    g392(.A(G2090), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n811), .A2(new_n812), .ZN(new_n821));
  NAND2_X1  g396(.A1(G299), .A2(G16), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n752), .A2(G20), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT23), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G1956), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n827), .ZN(new_n828));
  AOI211_X1 g403(.A(new_n814), .B(new_n828), .C1(new_n790), .C2(new_n789), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n781), .A2(new_n786), .A3(new_n792), .A4(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G6), .B(G305), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT32), .B(G1981), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT33), .B(G1976), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n530), .B1(new_n571), .B2(new_n602), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n608), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n606), .A2(new_n838), .A3(new_n607), .A4(new_n608), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n752), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n752), .B2(G23), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n833), .A2(KEYINPUT91), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(KEYINPUT91), .B2(new_n833), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n752), .A2(G22), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G166), .B2(new_n752), .ZN(new_n846));
  INV_X1    g421(.A(G1971), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n842), .B2(new_n834), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n844), .A2(KEYINPUT34), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n734), .A2(G25), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n495), .A2(G131), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n500), .A2(G119), .ZN(new_n853));
  OR2_X1    g428(.A1(G95), .A2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(G2104), .C1(G107), .C2(new_n480), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n851), .B1(new_n857), .B2(new_n734), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT89), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G1991), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  MUX2_X1   g436(.A(G24), .B(G290), .S(G16), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT90), .B(G1986), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n850), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT34), .B1(new_n844), .B2(new_n849), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(KEYINPUT36), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT36), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n830), .B1(new_n872), .B2(new_n873), .ZN(G311));
  INV_X1    g449(.A(new_n830), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n871), .B2(new_n876), .ZN(G150));
  NAND2_X1  g452(.A1(G80), .A2(G543), .ZN(new_n878));
  INV_X1    g453(.A(G67), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n571), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n880), .A2(new_n534), .B1(G93), .B2(new_n540), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n560), .A2(G55), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G860), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n652), .A2(G559), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT38), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n581), .A2(new_n881), .A3(new_n582), .A4(new_n882), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n582), .A2(new_n581), .B1(new_n881), .B2(new_n882), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n887), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT103), .ZN(new_n896));
  INV_X1    g471(.A(G860), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n885), .B1(new_n896), .B2(new_n898), .ZN(G145));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n497), .B(new_n677), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n504), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n510), .A2(new_n520), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n802), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n742), .A2(new_n772), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n774), .B2(new_n742), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n904), .B(new_n906), .C1(new_n774), .C2(new_n742), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n495), .A2(G142), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n500), .A2(G130), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n480), .A2(G118), .ZN(new_n912));
  OAI21_X1  g487(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n666), .B(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n856), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n909), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n908), .B2(new_n909), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n902), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n901), .B(G162), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n902), .A2(KEYINPUT105), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n917), .B1(new_n919), .B2(KEYINPUT104), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n908), .A2(new_n909), .A3(new_n927), .A4(new_n916), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n900), .B(new_n920), .C1(new_n925), .C2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(G166), .B(G305), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n837), .A2(new_n839), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n631), .A2(new_n636), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT79), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n623), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n840), .A2(new_n624), .A3(new_n631), .A4(new_n636), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(KEYINPUT107), .A3(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n935), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT108), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n940), .A2(KEYINPUT107), .A3(new_n941), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT107), .B1(new_n940), .B2(new_n941), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n947), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n933), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n650), .A2(G299), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n650), .A2(G299), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n650), .A2(G299), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT41), .B1(new_n961), .B2(new_n956), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n662), .A2(new_n892), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n891), .B1(new_n661), .B2(G559), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(new_n956), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT42), .B1(new_n952), .B2(new_n947), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n955), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n964), .A3(new_n965), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n967), .B2(new_n963), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n952), .A2(new_n953), .A3(new_n947), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n953), .B1(new_n952), .B2(new_n947), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT42), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n972), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(G868), .B1(new_n973), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n883), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G868), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n932), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n971), .B1(new_n955), .B2(new_n972), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n978), .A2(new_n975), .A3(new_n979), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n638), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n988), .A2(KEYINPUT109), .A3(new_n983), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n985), .A2(new_n989), .ZN(G295));
  NAND2_X1  g565(.A1(new_n981), .A2(new_n984), .ZN(G331));
  INV_X1    g566(.A(new_n968), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT110), .B1(new_n574), .B2(new_n575), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n574), .A2(KEYINPUT110), .A3(new_n575), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n994), .B(new_n995), .C1(new_n889), .C2(new_n890), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n583), .A2(new_n883), .ZN(new_n997));
  INV_X1    g572(.A(new_n995), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n888), .C1(new_n998), .C2(new_n993), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n996), .A2(G168), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G168), .B1(new_n996), .B2(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n992), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n999), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G286), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n999), .A3(G168), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n963), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(KEYINPUT111), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n963), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n976), .A2(new_n977), .ZN(new_n1012));
  AOI21_X1  g587(.A(G37), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n949), .A2(new_n954), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1006), .B(KEYINPUT112), .C1(new_n1008), .C2(new_n970), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1014), .B(new_n1015), .C1(KEYINPUT112), .C2(new_n1006), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1013), .A2(KEYINPUT43), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT43), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1013), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(G397));
  OR2_X1    g601(.A1(G290), .A2(G1986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(KEYINPUT113), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G137), .ZN(new_n1030));
  OAI221_X1 g605(.A(G40), .B1(new_n490), .B2(new_n491), .C1(new_n764), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n479), .B2(new_n484), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n522), .A2(new_n525), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1029), .B(new_n1040), .C1(KEYINPUT113), .C2(new_n1028), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT114), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1039), .B(KEYINPUT115), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n802), .A2(G2067), .ZN(new_n1044));
  INV_X1    g619(.A(G2067), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n797), .A2(new_n1045), .A3(new_n801), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n778), .B2(new_n772), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1039), .A2(G1996), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1043), .A2(new_n1048), .B1(new_n774), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n856), .B(new_n860), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1051), .B(KEYINPUT116), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1042), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1031), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1036), .A2(G1384), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1033), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n482), .A2(new_n483), .ZN(new_n1059));
  AOI211_X1 g634(.A(KEYINPUT67), .B(new_n480), .C1(new_n481), .C2(new_n476), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1056), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1384), .B1(new_n521), .B2(new_n527), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(KEYINPUT45), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n847), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n521), .A2(new_n527), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1034), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT50), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1035), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT117), .B(G2090), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1032), .A2(new_n1067), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G303), .A2(G8), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT55), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(G8), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1056), .B(new_n1068), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n840), .A2(G1976), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(G8), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT118), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1078), .A2(new_n1082), .A3(G8), .A4(new_n1079), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(KEYINPUT52), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n613), .A2(new_n617), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n613), .B2(new_n617), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1089), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1087), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1078), .A2(new_n1090), .A3(new_n1092), .A4(G8), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1078), .A2(G8), .A3(new_n1095), .A4(new_n1079), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1077), .A2(new_n1084), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1032), .A2(new_n1100), .A3(new_n1101), .A4(new_n1071), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1064), .B2(new_n1102), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1103), .A2(KEYINPUT119), .A3(new_n1076), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1076), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1066), .A2(new_n1036), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1032), .A2(new_n1108), .A3(new_n760), .A4(new_n1058), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1032), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n807), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1031), .A2(new_n1110), .A3(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(new_n1037), .A3(new_n478), .A4(new_n1058), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1109), .A2(new_n1110), .B1(new_n1112), .B2(new_n807), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1065), .A2(new_n1057), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1032), .A2(KEYINPUT53), .A3(new_n760), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(G301), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1107), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1116), .A2(G171), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(G301), .A3(new_n1120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1124), .A3(KEYINPUT54), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1070), .B1(new_n1069), .B2(new_n1062), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n790), .B(new_n1056), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1966), .B1(new_n1032), .B2(new_n1119), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G168), .A2(new_n1099), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1057), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1037), .B1(G164), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n751), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1032), .A2(new_n1067), .A3(new_n790), .A4(new_n1070), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(G8), .B(new_n1134), .C1(new_n1142), .C2(G286), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1131), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1136), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1106), .A2(new_n1122), .A3(new_n1125), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1112), .A2(new_n785), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1078), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1045), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT60), .ZN(new_n1151));
  INV_X1    g726(.A(new_n650), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT60), .A4(new_n650), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1150), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1032), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n826), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT56), .B(G2072), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1032), .A2(new_n1108), .A3(new_n1058), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n1162));
  OAI21_X1  g737(.A(G299), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1160), .A2(KEYINPUT123), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1157), .A2(new_n1165), .A3(new_n1159), .A4(KEYINPUT123), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1155), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1032), .A2(new_n1108), .A3(new_n778), .A4(new_n1058), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  XOR2_X1   g747(.A(KEYINPUT58), .B(G1341), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1078), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n584), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT59), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1167), .A2(KEYINPUT61), .A3(new_n1168), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1170), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1160), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1165), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1165), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n650), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1146), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1145), .A2(KEYINPUT62), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1136), .A2(new_n1143), .A3(new_n1188), .A4(new_n1144), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1106), .A2(new_n1187), .A3(new_n1121), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(G288), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1093), .A2(new_n1094), .A3(new_n1191), .ZN(new_n1192));
  AOI211_X1 g767(.A(new_n1099), .B(new_n1148), .C1(new_n1192), .C2(new_n1087), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1084), .A2(new_n1097), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1077), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1130), .A2(G286), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1106), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(KEYINPUT63), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1076), .B1(new_n1073), .B2(G8), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1200), .A2(new_n1098), .A3(new_n1201), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1190), .B(new_n1196), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1055), .B1(new_n1186), .B2(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1054), .A2(KEYINPUT127), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1054), .A2(KEYINPUT127), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1027), .A2(new_n1039), .ZN(new_n1207));
  XOR2_X1   g782(.A(new_n1207), .B(KEYINPUT48), .Z(new_n1208));
  NAND3_X1  g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1049), .B(KEYINPUT46), .Z(new_n1210));
  NAND2_X1  g785(.A1(new_n1047), .A2(new_n772), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1043), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT47), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n857), .A2(new_n860), .ZN(new_n1215));
  XOR2_X1   g790(.A(new_n1215), .B(KEYINPUT126), .Z(new_n1216));
  NAND2_X1  g791(.A1(new_n1050), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1046), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1043), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1209), .A2(new_n1214), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1204), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g796(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n929), .B1(new_n923), .B2(new_n924), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n920), .A2(new_n900), .ZN(new_n1225));
  OAI211_X1 g799(.A(new_n1223), .B(new_n697), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1227), .A2(KEYINPUT43), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1013), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(G308));
  NAND2_X1  g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  NAND4_X1  g805(.A1(new_n1231), .A2(new_n697), .A3(new_n930), .A4(new_n1223), .ZN(G225));
endmodule


