//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT69), .B(G238), .Z(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT68), .B(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n219), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n210), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n215), .B1(new_n216), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n216), .B2(new_n230), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  INV_X1    g0036(.A(G50), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n204), .A2(new_n205), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n237), .B1(new_n238), .B2(KEYINPUT66), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n239), .B1(KEYINPUT66), .B2(new_n238), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT67), .Z(new_n241));
  AOI21_X1  g0041(.A(new_n232), .B1(new_n236), .B2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n225), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n237), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n202), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT70), .B1(new_n258), .B2(new_n233), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT70), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G1), .A4(G13), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G226), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G222), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G223), .A2(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n258), .A2(new_n233), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n272), .B(new_n273), .C1(G77), .C2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(new_n264), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n259), .A2(new_n275), .A3(G274), .A4(new_n262), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n265), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT71), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(new_n233), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n208), .A2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n289), .B1(G50), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  XOR2_X1   g0091(.A(KEYINPUT8), .B(G58), .Z(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n209), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n209), .B1(new_n238), .B2(new_n237), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(KEYINPUT72), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n302), .B2(new_n285), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n283), .B(new_n303), .C1(G179), .C2(new_n281), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n279), .B2(new_n280), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G200), .B2(new_n281), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n303), .B(KEYINPUT9), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n284), .A2(new_n233), .ZN(new_n313));
  INV_X1    g0113(.A(new_n218), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n209), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n297), .A2(new_n237), .B1(new_n294), .B2(new_n226), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  INV_X1    g0120(.A(new_n287), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G68), .A3(new_n288), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n314), .B2(new_n286), .ZN(new_n324));
  OR2_X1    g0124(.A1(KEYINPUT12), .A2(G68), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n286), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n319), .A2(new_n320), .A3(new_n322), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n234), .A2(new_n260), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n268), .A2(KEYINPUT74), .A3(G226), .A4(new_n269), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT74), .ZN(new_n335));
  AND2_X1   g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  NOR2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n269), .A2(G226), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n329), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n263), .A2(G238), .A3(new_n264), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n276), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT13), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n328), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n342), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n345), .A3(G179), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n345), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n328), .B1(new_n355), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n327), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n327), .B1(new_n355), .B2(G200), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n305), .B2(new_n355), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n217), .A2(new_n269), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n268), .B1(new_n225), .B2(G1698), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n273), .B1(G107), .B2(new_n268), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n263), .A2(G244), .A3(new_n264), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n276), .A3(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(G179), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n282), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n293), .A2(new_n297), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n368), .A2(new_n294), .B1(new_n209), .B2(new_n226), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n313), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n226), .B1(new_n208), .B2(G20), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n286), .A2(KEYINPUT73), .A3(G77), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT73), .B1(new_n286), .B2(G77), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n321), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n364), .A2(G200), .ZN(new_n377));
  INV_X1    g0177(.A(new_n375), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n305), .C2(new_n364), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n357), .A2(new_n359), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n292), .A2(new_n288), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(new_n287), .B1(new_n286), .B2(new_n292), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT77), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n259), .A2(G232), .A3(new_n264), .A4(new_n262), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(G1698), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n268), .B1(G33), .B2(G87), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n276), .B(new_n386), .C1(new_n390), .C2(new_n329), .ZN(new_n391));
  INV_X1    g0191(.A(G200), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(G1698), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G223), .B2(G1698), .ZN(new_n395));
  INV_X1    g0195(.A(G33), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n395), .A2(new_n338), .B1(new_n396), .B2(new_n221), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n273), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n398), .A2(new_n305), .A3(new_n276), .A4(new_n386), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n204), .B(new_n205), .C1(new_n218), .C2(new_n202), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(G20), .B1(G159), .B2(new_n296), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n338), .B2(new_n209), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n267), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n313), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n338), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n266), .A2(new_n209), .A3(new_n267), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n314), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT16), .B1(new_n416), .B2(new_n402), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n385), .B(new_n400), .C1(new_n408), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n203), .A2(KEYINPUT68), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT68), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n202), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n423), .B2(new_n238), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n296), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n314), .B2(new_n415), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n313), .B(new_n407), .C1(new_n427), .C2(KEYINPUT16), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n385), .A4(new_n400), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n385), .B1(new_n408), .B2(new_n417), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n391), .A2(G169), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n398), .A2(G179), .A3(new_n276), .A4(new_n386), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT18), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n435), .B1(new_n428), .B2(new_n385), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n431), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n312), .A2(new_n382), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G283), .ZN(new_n444));
  AND2_X1   g0244(.A1(KEYINPUT78), .A2(G97), .ZN(new_n445));
  NOR2_X1   g0245(.A1(KEYINPUT78), .A2(G97), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n209), .B(new_n444), .C1(new_n447), .C2(G33), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT20), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  AOI22_X1  g0250(.A1(KEYINPUT82), .A2(new_n449), .B1(new_n450), .B2(G20), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n449), .A2(KEYINPUT82), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n448), .A2(new_n313), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n286), .A2(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n208), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n286), .A2(new_n456), .A3(new_n233), .A4(new_n284), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n450), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n444), .A2(new_n209), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT78), .B(G97), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n396), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(new_n313), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n452), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n454), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G41), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n208), .B(G45), .C1(new_n466), .C2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(G274), .A3(new_n259), .A4(new_n262), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n269), .A2(G257), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G264), .A2(G1698), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n336), .C2(new_n337), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(new_n273), .C1(G303), .C2(new_n268), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n468), .A2(G41), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n208), .A4(G45), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(new_n259), .A3(G270), .A4(new_n262), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n471), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n465), .A2(KEYINPUT21), .A3(G169), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT83), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(G169), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT21), .A4(new_n465), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n465), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n487), .A2(new_n488), .B1(new_n465), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n465), .B1(G200), .B2(new_n480), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n305), .B2(new_n480), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(new_n269), .C1(new_n336), .C2(new_n337), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n268), .A2(KEYINPUT86), .A3(G250), .A4(new_n269), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(G1698), .C1(new_n336), .C2(new_n337), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G294), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n329), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n478), .A2(new_n259), .A3(G264), .A4(new_n262), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n471), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n489), .ZN(new_n508));
  INV_X1    g0308(.A(new_n506), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n502), .B1(new_n497), .B2(new_n498), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n329), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n282), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n209), .B(G87), .C1(new_n336), .C2(new_n337), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n268), .A2(new_n516), .A3(new_n209), .A4(G87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT84), .B1(new_n520), .B2(G20), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n520), .A2(KEYINPUT84), .A3(G20), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n513), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n525), .A3(new_n513), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n285), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n286), .ZN(new_n530));
  INV_X1    g0330(.A(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n536), .B1(G107), .B2(new_n458), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n508), .B(new_n512), .C1(new_n529), .C2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n518), .A2(new_n525), .A3(new_n513), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n313), .B1(new_n540), .B2(new_n526), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n509), .B(G190), .C1(new_n510), .C2(new_n329), .ZN(new_n542));
  OAI21_X1  g0342(.A(G200), .B1(new_n504), .B2(new_n506), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n537), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n209), .B1(new_n331), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(KEYINPUT78), .A2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT78), .A2(G97), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n531), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g0350(.A(KEYINPUT80), .B(G87), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n268), .A2(new_n209), .A3(G68), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n546), .B1(new_n447), .B2(new_n294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT81), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n552), .A2(new_n554), .A3(new_n557), .A4(new_n553), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n313), .A3(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n457), .A2(new_n368), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n368), .A2(new_n530), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G45), .ZN(new_n563));
  OR3_X1    g0363(.A1(new_n563), .A2(G1), .A3(G274), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n222), .B1(new_n563), .B2(G1), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n259), .A2(new_n564), .A3(new_n262), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(G238), .A2(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n227), .A2(G1698), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n336), .C2(new_n337), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n329), .B1(new_n570), .B2(new_n520), .ZN(new_n571));
  OAI21_X1  g0371(.A(G169), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G238), .A2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n227), .B2(G1698), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n268), .B1(G33), .B2(G116), .ZN(new_n575));
  OAI211_X1 g0375(.A(G179), .B(new_n566), .C1(new_n575), .C2(new_n329), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n562), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n566), .B1(new_n575), .B2(new_n329), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n392), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n579), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n458), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n561), .A3(new_n559), .A4(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n227), .A2(G1698), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n336), .B2(new_n337), .ZN(new_n586));
  NOR2_X1   g0386(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(new_n587), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n590), .B(new_n585), .C1(new_n337), .C2(new_n336), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n444), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n273), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n478), .A2(new_n259), .A3(G257), .A4(new_n262), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n471), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n415), .A2(G107), .ZN(new_n598));
  XOR2_X1   g0398(.A(G97), .B(G107), .Z(new_n599));
  NAND2_X1  g0399(.A1(new_n531), .A2(KEYINPUT6), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(KEYINPUT6), .B1(new_n447), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n313), .ZN(new_n604));
  INV_X1    g0404(.A(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n530), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n457), .B2(new_n605), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n593), .A2(new_n595), .A3(G190), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n597), .A2(new_n604), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n593), .A2(new_n595), .A3(G179), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n282), .B1(new_n593), .B2(new_n595), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n285), .B1(new_n598), .B2(new_n602), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(new_n607), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n584), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n443), .A2(new_n494), .A3(new_n545), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n304), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n359), .A2(new_n366), .A3(new_n365), .A4(new_n375), .ZN(new_n619));
  INV_X1    g0419(.A(new_n357), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n431), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n438), .A3(new_n441), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n310), .A2(new_n311), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n559), .A2(new_n561), .A3(new_n582), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n572), .A2(KEYINPUT87), .A3(new_n576), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT87), .B1(new_n572), .B2(new_n576), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n625), .A2(new_n581), .B1(new_n628), .B2(new_n562), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n613), .A2(new_n607), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT88), .B1(new_n611), .B2(new_n612), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n596), .A2(G169), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT88), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n593), .A2(new_n595), .A3(G179), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n630), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n629), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n634), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n578), .A2(new_n639), .A3(new_n583), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n628), .A2(new_n562), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n638), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT89), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT89), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n638), .A2(new_n646), .A3(new_n642), .A4(new_n643), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n610), .A2(new_n544), .A3(new_n614), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n629), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n539), .A2(new_n486), .A3(new_n491), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n645), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n443), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n624), .A2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n465), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n494), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n486), .A2(new_n491), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n662), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n661), .B1(new_n529), .B2(new_n538), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n545), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n661), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n539), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n666), .A2(KEYINPUT90), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n539), .A2(new_n661), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n664), .A2(new_n661), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n545), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n212), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G1), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n550), .A2(new_n551), .A3(G116), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n240), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n629), .A2(new_n636), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(new_n614), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n584), .A2(new_n637), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n689), .A3(new_n643), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT91), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n664), .A2(new_n691), .A3(new_n539), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n651), .A2(KEYINPUT91), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n649), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT29), .B(new_n669), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n644), .A2(KEYINPUT89), .B1(new_n650), .B2(new_n651), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n661), .B1(new_n696), .B2(new_n647), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n695), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n616), .A2(new_n494), .A3(new_n545), .A4(new_n669), .ZN(new_n699));
  INV_X1    g0499(.A(new_n596), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n475), .A2(new_n479), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n576), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n507), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n700), .A2(KEYINPUT30), .A3(new_n507), .A4(new_n702), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n579), .A2(new_n489), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n511), .A2(new_n596), .A3(new_n480), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n661), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n699), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n698), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n685), .B1(new_n718), .B2(G1), .ZN(G364));
  NOR2_X1   g0519(.A1(new_n211), .A2(G20), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n208), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n680), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n212), .A2(new_n338), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G355), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G116), .B2(new_n213), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n241), .A2(new_n563), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n212), .A2(new_n268), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n253), .B2(G45), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n209), .B1(KEYINPUT92), .B2(new_n282), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n282), .A2(KEYINPUT92), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n233), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n723), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(G20), .A2(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT93), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n209), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT94), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G326), .A2(new_n749), .B1(new_n756), .B2(G303), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n742), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n268), .B1(new_n760), .B2(G311), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n750), .A2(new_n758), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n741), .A2(new_n305), .A3(G200), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n763), .A2(G329), .B1(new_n764), .B2(G322), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n741), .A2(new_n392), .A3(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(KEYINPUT33), .B(G317), .Z(new_n768));
  NAND3_X1  g0568(.A1(new_n750), .A2(new_n305), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n209), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(G294), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n757), .A2(new_n761), .A3(new_n765), .A4(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n760), .A2(G77), .B1(G58), .B2(new_n764), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n605), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n763), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G68), .C2(new_n766), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n237), .B2(new_n748), .ZN(new_n782));
  INV_X1    g0582(.A(new_n769), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G107), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n268), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n756), .B2(new_n551), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT95), .Z(new_n787));
  OAI21_X1  g0587(.A(new_n776), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n740), .B1(new_n788), .B2(new_n734), .ZN(new_n789));
  INV_X1    g0589(.A(new_n737), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n665), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n666), .ZN(new_n792));
  INV_X1    g0592(.A(new_n723), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n665), .A2(G330), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(G396));
  NAND3_X1  g0596(.A1(new_n653), .A2(new_n381), .A3(new_n669), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n379), .B1(new_n378), .B2(new_n669), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n376), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n376), .A2(new_n661), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n797), .B1(new_n697), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(new_n716), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n723), .B1(new_n802), .B2(new_n716), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n734), .A2(new_n735), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n793), .B1(new_n806), .B2(new_n226), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n801), .A2(new_n736), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n769), .A2(new_n221), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G311), .A2(new_n763), .B1(new_n760), .B2(G116), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n770), .B2(new_n767), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n810), .B(new_n812), .C1(G303), .C2(new_n749), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n268), .B1(new_n756), .B2(G107), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT96), .ZN(new_n815));
  INV_X1    g0615(.A(new_n764), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n773), .A2(new_n605), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n813), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n814), .A2(KEYINPUT96), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n268), .B1(new_n762), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT100), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n773), .A2(new_n202), .B1(new_n769), .B2(new_n203), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT98), .B(G143), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n760), .A2(G159), .B1(new_n828), .B2(new_n764), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n295), .B2(new_n767), .C1(new_n748), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n826), .B1(new_n237), .B2(new_n755), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n831), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n832), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n820), .A2(new_n821), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n808), .B(new_n809), .C1(new_n734), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n805), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  OR2_X1    g0640(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(G116), .A3(new_n236), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  OAI21_X1  g0644(.A(G77), .B1(new_n218), .B2(new_n202), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n240), .A2(new_n845), .B1(G50), .B2(new_n203), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n208), .A2(G13), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G330), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n327), .A2(new_n661), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n357), .A2(new_n359), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n327), .B(new_n661), .C1(new_n354), .C2(new_n356), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n714), .A2(new_n853), .A3(new_n801), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n659), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n432), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n442), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n437), .A2(new_n857), .A3(new_n861), .A4(new_n418), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n418), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT102), .B1(new_n864), .B2(new_n439), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n437), .A2(new_n866), .A3(new_n418), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n869), .B2(KEYINPUT103), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n437), .A2(new_n418), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n858), .B1(new_n871), .B2(KEYINPUT102), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n861), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n860), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(new_n408), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n402), .A2(new_n406), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(KEYINPUT16), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n880), .A2(new_n385), .B1(new_n435), .B2(new_n659), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n881), .B2(new_n864), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n862), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n659), .B1(new_n880), .B2(new_n385), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n442), .A2(KEYINPUT101), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT101), .B1(new_n442), .B2(new_n884), .ZN(new_n886));
  OAI211_X1 g0686(.A(KEYINPUT38), .B(new_n883), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT40), .B(new_n855), .C1(new_n877), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n854), .B1(new_n892), .B2(new_n887), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n889), .B1(KEYINPUT40), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n443), .A2(new_n714), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT104), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n849), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n620), .A2(new_n669), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n887), .C1(new_n876), .C2(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n442), .A2(new_n884), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT101), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n442), .A2(KEYINPUT101), .A3(new_n884), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n907), .B2(new_n883), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT39), .B1(new_n908), .B2(new_n888), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n900), .B1(new_n902), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n853), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n797), .B2(new_n800), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n892), .A2(new_n887), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n438), .A2(new_n441), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n914), .B1(new_n915), .B2(new_n659), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n443), .B(new_n695), .C1(new_n697), .C2(KEYINPUT29), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n624), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n899), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n208), .B2(new_n720), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n899), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n848), .B1(new_n922), .B2(new_n923), .ZN(G367));
  AND2_X1   g0724(.A1(new_n249), .A2(new_n728), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n738), .B1(new_n213), .B2(new_n368), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n723), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n767), .A2(new_n817), .B1(new_n769), .B2(new_n447), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n268), .B1(G303), .B2(new_n764), .ZN(new_n929));
  INV_X1    g0729(.A(G317), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n929), .B1(new_n770), .B2(new_n759), .C1(new_n930), .C2(new_n762), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n928), .B(new_n931), .C1(G107), .C2(new_n774), .ZN(new_n932));
  INV_X1    g0732(.A(G311), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n933), .B2(new_n748), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n755), .A2(new_n450), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT46), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n774), .A2(G68), .B1(new_n764), .B2(G150), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n748), .B2(new_n827), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT107), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n268), .B1(new_n762), .B2(new_n830), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n760), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n783), .A2(G77), .B1(new_n766), .B2(G159), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n755), .C2(new_n202), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n934), .A2(new_n936), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n927), .B1(new_n945), .B2(new_n734), .ZN(new_n946));
  INV_X1    g0746(.A(new_n643), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n625), .A2(new_n669), .ZN(new_n948));
  MUX2_X1   g0748(.A(new_n629), .B(new_n947), .S(new_n948), .Z(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n790), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n673), .A2(new_n674), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n615), .B1(new_n630), .B2(new_n669), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n636), .A2(new_n661), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n678), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n678), .A2(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n675), .A2(new_n959), .A3(new_n956), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n677), .A2(new_n545), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n670), .B2(new_n677), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n666), .B(new_n965), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n718), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n680), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n722), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n952), .A2(new_n953), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n539), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n669), .B1(new_n972), .B2(new_n688), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n971), .B2(new_n964), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n954), .A2(new_n545), .A3(new_n677), .A4(new_n974), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(KEYINPUT106), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n949), .B(KEYINPUT43), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n982), .A2(new_n984), .B1(new_n675), .B2(new_n971), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n675), .A2(new_n971), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n979), .A2(new_n981), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n983), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n950), .B1(new_n970), .B2(new_n990), .ZN(G387));
  AOI21_X1  g0791(.A(new_n729), .B1(new_n246), .B2(G45), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n683), .B2(new_n724), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n292), .A2(new_n237), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT50), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n563), .B1(new_n203), .B2(new_n226), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n995), .A2(new_n683), .A3(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n993), .A2(new_n997), .B1(G107), .B2(new_n213), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n793), .B1(new_n998), .B2(new_n738), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n773), .A2(new_n368), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n293), .B2(new_n767), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G97), .B2(new_n783), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n762), .A2(new_n295), .B1(new_n759), .B2(new_n203), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n338), .B(new_n1004), .C1(G50), .C2(new_n764), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n749), .A2(G159), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n756), .A2(G77), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n268), .B1(new_n763), .B2(G326), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n755), .A2(new_n817), .B1(new_n770), .B2(new_n773), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n760), .A2(G303), .B1(G317), .B2(new_n764), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n933), .B2(new_n767), .C1(new_n748), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1009), .B1(new_n450), .B2(new_n769), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1008), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n734), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n999), .B(new_n1021), .C1(new_n670), .C2(new_n790), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT108), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n966), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n718), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n680), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n718), .A2(new_n1024), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1023), .B1(new_n721), .B2(new_n966), .C1(new_n1026), .C2(new_n1027), .ZN(G393));
  AOI22_X1  g0828(.A1(new_n749), .A2(G150), .B1(G159), .B2(new_n764), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT110), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT51), .Z(new_n1031));
  NOR2_X1   g0831(.A1(new_n755), .A2(new_n218), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n268), .B1(new_n762), .B2(new_n827), .C1(new_n293), .C2(new_n759), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n810), .B1(G50), .B2(new_n766), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n226), .B2(new_n773), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT111), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n748), .A2(new_n930), .B1(new_n933), .B2(new_n816), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n338), .B1(new_n759), .B2(new_n817), .C1(new_n1012), .C2(new_n762), .ZN(new_n1040));
  INV_X1    g0840(.A(G303), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n784), .B1(new_n1041), .B2(new_n767), .C1(new_n450), .C2(new_n773), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(G283), .C2(new_n756), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT112), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n734), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n971), .A2(new_n737), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n739), .B1(new_n212), .B2(new_n461), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n256), .A2(new_n728), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n793), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT109), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n961), .A2(new_n962), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n951), .A2(new_n960), .A3(KEYINPUT109), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1055), .B2(new_n722), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1053), .A2(new_n1025), .A3(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n680), .B1(new_n963), .B2(new_n1025), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n851), .A2(new_n1060), .A3(new_n852), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n851), .B2(new_n852), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n714), .A2(G330), .A3(new_n801), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n669), .B(new_n799), .C1(new_n690), .C2(new_n694), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n715), .A2(new_n801), .A3(new_n853), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1065), .A2(new_n800), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1064), .A2(new_n912), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n797), .A2(new_n800), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n715), .A2(new_n443), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n624), .A2(new_n918), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n900), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n902), .B(new_n909), .C1(new_n913), .C2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1066), .A2(new_n800), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n888), .B2(new_n877), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1079), .A2(new_n1083), .A3(new_n1067), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1067), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1067), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1075), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1079), .A2(new_n1083), .A3(new_n1067), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1086), .A2(new_n1092), .A3(new_n680), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n722), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n774), .A2(G159), .B1(new_n766), .B2(G137), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(KEYINPUT54), .B(G143), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT114), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1099), .B2(new_n759), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT115), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n755), .A2(new_n295), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n338), .B1(new_n763), .B2(G125), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n237), .B2(new_n769), .C1(new_n822), .C2(new_n816), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G128), .B2(new_n749), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n760), .A2(new_n461), .B1(G107), .B2(new_n766), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n748), .B2(new_n770), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n338), .B1(new_n755), .B2(new_n221), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n773), .A2(new_n226), .B1(new_n816), .B2(new_n450), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT118), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n769), .A2(new_n203), .B1(new_n762), .B2(new_n817), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n734), .B1(new_n1108), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n793), .B1(new_n806), .B2(new_n293), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n902), .A2(new_n909), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1119), .C1(new_n1120), .C2(new_n736), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1093), .A2(new_n1095), .A3(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n913), .A2(new_n914), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n915), .A2(new_n659), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n910), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n914), .A2(new_n855), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT40), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n849), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n623), .A2(new_n304), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n303), .A2(new_n856), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n312), .A2(new_n1130), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1129), .A2(new_n889), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(G330), .B1(new_n893), .B2(KEYINPUT40), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n714), .A2(new_n853), .A3(KEYINPUT40), .A4(new_n801), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n862), .B1(new_n873), .B2(new_n874), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n869), .A2(KEYINPUT103), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n859), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n891), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n1146), .B2(new_n887), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1138), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1126), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1140), .A2(new_n1148), .B1(new_n911), .B2(new_n916), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT57), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1075), .B1(new_n1094), .B2(new_n1073), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n680), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1092), .A2(new_n1076), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1139), .B1(new_n1129), .B2(new_n889), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1141), .A2(new_n1147), .A3(new_n1138), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n917), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1126), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1153), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n735), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n268), .A2(G41), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n237), .B1(G33), .B2(G41), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n748), .A2(new_n450), .B1(new_n203), .B2(new_n773), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n767), .A2(new_n605), .B1(new_n368), .B2(new_n759), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT119), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1163), .B1(new_n770), .B2(new_n762), .C1(new_n531), .C2(new_n816), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G58), .B2(new_n783), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1167), .A2(new_n1007), .A3(new_n1169), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n760), .A2(G137), .B1(G128), .B2(new_n764), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n822), .B2(new_n767), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G150), .B2(new_n774), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n749), .A2(G125), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n755), .C2(new_n1099), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n783), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1174), .B1(new_n1173), .B2(new_n1172), .C1(new_n1180), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n734), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT121), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n793), .B(new_n1187), .C1(new_n237), .C2(new_n806), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1159), .A2(new_n722), .B1(new_n1162), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1161), .A2(new_n1189), .ZN(G375));
  AOI21_X1  g0990(.A(new_n793), .B1(new_n806), .B2(new_n203), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n338), .B1(new_n759), .B2(new_n531), .C1(new_n816), .C2(new_n770), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1001), .B1(new_n226), .B2(new_n769), .C1(new_n450), .C2(new_n767), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G294), .C2(new_n749), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n755), .A2(new_n605), .B1(new_n1041), .B2(new_n762), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT122), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n773), .A2(new_n237), .B1(new_n769), .B2(new_n202), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n763), .A2(G128), .B1(new_n764), .B2(G137), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n268), .C1(new_n295), .C2(new_n759), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n766), .C2(new_n1098), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G132), .A2(new_n749), .B1(new_n756), .B2(G159), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1194), .A2(new_n1196), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n734), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1191), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1063), .B2(new_n735), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1073), .B2(new_n722), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1077), .A2(new_n969), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT123), .Z(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G381));
  NOR3_X1   g1011(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n970), .A2(new_n990), .ZN(new_n1214));
  INV_X1    g1014(.A(G390), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n950), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G378), .A2(G375), .A3(new_n1213), .A4(new_n1216), .ZN(G407));
  INV_X1    g1017(.A(G213), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(G343), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(G375), .A2(G378), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT124), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1023(.A(G378), .B(new_n1189), .C1(new_n1153), .C2(new_n1160), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n968), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT125), .B1(new_n1226), .B2(new_n1154), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n722), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1188), .A2(new_n1162), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1154), .A3(KEYINPUT125), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G378), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1220), .B1(new_n1225), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1208), .A2(KEYINPUT60), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT60), .A4(new_n1075), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1077), .A2(new_n680), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1206), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1219), .A2(G2897), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1238), .B(new_n839), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT61), .B1(new_n1234), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n969), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1152), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1189), .A3(new_n1232), .ZN(new_n1250));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1219), .B1(new_n1252), .B2(new_n1224), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1239), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1220), .B(new_n1239), .C1(new_n1225), .C2(new_n1233), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1246), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(G393), .B(G396), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(G390), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1216), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1216), .B2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT127), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1263), .B(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1263), .B(new_n1267), .C1(new_n1253), .C2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1219), .B(new_n1242), .C1(new_n1252), .C2(new_n1224), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1272), .B2(KEYINPUT63), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(KEYINPUT63), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1256), .A2(KEYINPUT126), .A3(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1270), .A2(new_n1273), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1266), .A2(new_n1277), .ZN(G405));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1251), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1224), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1239), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1224), .A3(new_n1242), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1263), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1263), .A3(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


