//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(new_n211), .B2(new_n212), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n218), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n247), .A2(new_n206), .A3(G1), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n213), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n205), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n206), .B1(new_n201), .B2(new_n249), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G20), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI211_X1 g0065(.A(new_n257), .B(new_n261), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n252), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n250), .B1(new_n254), .B2(new_n256), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  AND2_X1   g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G41), .A2(G45), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n270), .A2(new_n213), .B1(new_n271), .B2(G1), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT65), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT65), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  AND2_X1   g0087(.A1(G1), .A2(G13), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n275), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n289), .A3(new_n205), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n276), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G222), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(G1698), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n280), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n268), .A2(new_n269), .B1(G200), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n302), .B1(new_n269), .B2(new_n268), .C1(new_n303), .C2(new_n301), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT10), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n301), .A2(G179), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n268), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n291), .A2(new_n293), .ZN(new_n311));
  INV_X1    g0111(.A(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n298), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(G226), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G87), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n276), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n290), .B1(new_n232), .B2(new_n272), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  OR3_X1    g0121(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n265), .A2(new_n255), .ZN(new_n325));
  INV_X1    g0125(.A(new_n248), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n254), .A2(new_n325), .B1(new_n326), .B2(new_n265), .ZN(new_n327));
  INV_X1    g0127(.A(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n220), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n201), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n258), .A2(G159), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n311), .B2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n294), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n336), .B2(G68), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n267), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n293), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT7), .B(new_n206), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n220), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n344), .B2(new_n332), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n327), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT18), .B1(new_n324), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n327), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n334), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G68), .ZN(new_n350));
  INV_X1    g0150(.A(new_n332), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT16), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n335), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT7), .B1(new_n294), .B2(new_n206), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n351), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n252), .B1(new_n356), .B2(new_n339), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n348), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n323), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n347), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n317), .B2(new_n318), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n319), .B2(G190), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n348), .C1(new_n357), .C2(new_n352), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n346), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n253), .A2(G77), .A3(new_n255), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n264), .A2(new_n259), .B1(new_n206), .B2(new_n295), .ZN(new_n371));
  XOR2_X1   g0171(.A(KEYINPUT15), .B(G87), .Z(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n263), .B2(new_n372), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n370), .B1(G77), .B2(new_n326), .C1(new_n373), .C2(new_n267), .ZN(new_n374));
  INV_X1    g0174(.A(new_n276), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n294), .A2(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G232), .ZN(new_n377));
  INV_X1    g0177(.A(G107), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n311), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n294), .A2(new_n221), .A3(new_n312), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n279), .A2(G244), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n290), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n374), .B1(new_n384), .B2(G190), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n362), .B2(new_n384), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n307), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(new_n374), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n321), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n310), .A2(new_n361), .A3(new_n369), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n258), .A2(G50), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT68), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n263), .A2(G77), .B1(G20), .B2(new_n220), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n267), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(KEYINPUT11), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n326), .A2(KEYINPUT12), .A3(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT12), .B1(new_n326), .B2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n220), .B1(new_n205), .B2(G20), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n399), .A2(new_n400), .B1(new_n253), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n232), .A2(G1698), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n311), .B(new_n406), .C1(G226), .C2(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n276), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n221), .B1(new_n274), .B2(new_n278), .ZN(new_n411));
  INV_X1    g0211(.A(new_n290), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n411), .A2(KEYINPUT67), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT67), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n277), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT66), .B1(new_n276), .B2(new_n277), .ZN(new_n416));
  OAI21_X1  g0216(.A(G238), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n417), .B2(new_n290), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n410), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT67), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n417), .A2(new_n414), .A3(new_n290), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n410), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n307), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n405), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n423), .B2(new_n410), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT13), .B(new_n409), .C1(new_n421), .C2(new_n422), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT70), .A3(KEYINPUT14), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n420), .A2(G179), .A3(new_n425), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n420), .A2(new_n436), .A3(G179), .A4(new_n425), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n435), .A2(new_n437), .B1(new_n427), .B2(new_n426), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT72), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n433), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n433), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n404), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n429), .A2(new_n430), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G190), .ZN(new_n444));
  OAI21_X1  g0244(.A(G200), .B1(new_n429), .B2(new_n430), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n403), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT69), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT69), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n448), .A3(new_n403), .A4(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n392), .A2(new_n442), .A3(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n291), .A2(new_n293), .A3(new_n206), .A4(G87), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT22), .ZN(new_n453));
  XOR2_X1   g0253(.A(KEYINPUT80), .B(KEYINPUT24), .Z(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n206), .B2(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n378), .A2(KEYINPUT23), .A3(G20), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n453), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n455), .B1(new_n453), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n252), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n253), .B1(G1), .B2(new_n262), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT25), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n326), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n378), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n466), .A2(G107), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT81), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n464), .A2(KEYINPUT81), .A3(new_n470), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n311), .A2(G257), .A3(G1698), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n311), .A2(G250), .A3(new_n312), .ZN(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n262), .C2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n205), .B(G45), .C1(new_n478), .C2(G41), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n282), .A2(new_n284), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n478), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n375), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n477), .A2(new_n375), .B1(new_n482), .B2(G264), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n289), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G169), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n321), .B2(new_n485), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n472), .A2(new_n473), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(G200), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(G190), .A3(new_n484), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n464), .A3(new_n470), .A4(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n248), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n465), .B2(new_n493), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n349), .A2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n378), .A2(KEYINPUT6), .A3(G97), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n493), .A2(new_n378), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(G20), .B1(G77), .B2(new_n258), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n495), .B1(new_n503), .B2(new_n252), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n481), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G257), .A3(new_n276), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n507), .A2(new_n484), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n311), .A2(G250), .A3(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n311), .A2(G244), .A3(new_n312), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT4), .B1(new_n376), .B2(G244), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n375), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT75), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n508), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n505), .B1(new_n520), .B2(G190), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(KEYINPUT74), .B(new_n375), .C1(new_n513), .C2(new_n514), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n508), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n517), .A2(new_n307), .A3(new_n519), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n507), .A2(new_n484), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n523), .B2(new_n524), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n504), .B1(new_n530), .B2(new_n321), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n521), .A2(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n492), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n482), .A2(G270), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n484), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n311), .A2(G264), .A3(G1698), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n311), .A2(G257), .A3(new_n312), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n294), .A2(G303), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n276), .B1(new_n541), .B2(KEYINPUT79), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n535), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n510), .B(new_n206), .C1(G33), .C2(new_n493), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n252), .C1(new_n206), .C2(G116), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT20), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n248), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n465), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g0349(.A(G169), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT21), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n540), .ZN(new_n552));
  INV_X1    g0352(.A(new_n535), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n550), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT21), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n543), .B(G179), .C1(new_n546), .C2(new_n549), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n553), .A3(G190), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n546), .A2(new_n549), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n560), .B(new_n561), .C1(new_n543), .C2(new_n362), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n311), .A2(new_n206), .A3(G68), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n311), .A2(KEYINPUT76), .A3(new_n206), .A4(G68), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n263), .A2(new_n568), .A3(G97), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n499), .A2(new_n222), .B1(new_n408), .B2(new_n206), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n568), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n372), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n252), .B1(new_n248), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n466), .A2(new_n372), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n574), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n223), .B1(new_n285), .B2(G1), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n205), .A2(new_n287), .A3(G45), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n276), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n311), .A2(G238), .A3(new_n312), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n311), .A2(G244), .A3(G1698), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n456), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(new_n586), .B2(new_n375), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G179), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n307), .B2(new_n587), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n577), .A2(new_n579), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n572), .A2(new_n252), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n573), .A2(new_n248), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n466), .A2(G87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n362), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n587), .A2(G190), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n595), .A2(new_n596), .A3(new_n591), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n590), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n563), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n451), .A2(new_n533), .A3(new_n603), .ZN(G372));
  INV_X1    g0404(.A(KEYINPUT83), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n426), .A2(new_n405), .A3(new_n427), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT70), .B1(new_n431), .B2(KEYINPUT14), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n426), .A2(new_n427), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n436), .B1(new_n443), .B2(G179), .ZN(new_n610));
  INV_X1    g0410(.A(new_n437), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT72), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n433), .A2(new_n438), .A3(new_n439), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n403), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n390), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n446), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n605), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n365), .A2(new_n366), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT17), .B1(new_n346), .B2(new_n364), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n617), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n347), .A2(new_n360), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n305), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n309), .ZN(new_n628));
  INV_X1    g0428(.A(new_n451), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n464), .A2(new_n470), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n487), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(new_n558), .A3(new_n559), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT82), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n587), .A2(new_n307), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n321), .B(new_n583), .C1(new_n586), .C2(new_n375), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n588), .B(KEYINPUT82), .C1(new_n307), .C2(new_n587), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n576), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n595), .A2(new_n596), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n598), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(new_n491), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n532), .A2(new_n632), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n531), .A2(new_n638), .A3(new_n528), .A4(new_n640), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n531), .A2(new_n528), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT26), .B1(new_n601), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n642), .A2(new_n644), .A3(new_n646), .A4(new_n638), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n628), .A2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n558), .A2(new_n559), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(KEYINPUT84), .B(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n473), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n471), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n487), .A3(new_n656), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n656), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n492), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n661), .B1(new_n663), .B2(new_n660), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n650), .B(new_n657), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n631), .A2(new_n656), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n561), .A2(new_n657), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n563), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(G399));
  AND2_X1   g0478(.A1(new_n282), .A2(new_n284), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n209), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n499), .A2(new_n222), .A3(new_n547), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n215), .B2(new_n680), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n508), .A2(new_n515), .A3(new_n518), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n518), .B1(new_n508), .B2(new_n515), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n543), .A2(new_n483), .A3(new_n635), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n543), .A2(new_n483), .A3(new_n635), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n520), .A3(KEYINPUT30), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n587), .B(KEYINPUT86), .ZN(new_n695));
  AOI21_X1  g0495(.A(G179), .B1(new_n483), .B2(new_n484), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n526), .A2(new_n695), .A3(new_n554), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n692), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n656), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT87), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n602), .A2(new_n492), .A3(new_n532), .A4(new_n657), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT31), .B1(new_n698), .B2(new_n656), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT87), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n686), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n647), .A2(new_n657), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT88), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT88), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n647), .A2(new_n714), .A3(new_n657), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n601), .A2(new_n645), .A3(KEYINPUT26), .ZN(new_n717));
  INV_X1    g0517(.A(new_n638), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n532), .A2(new_n641), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n650), .B1(new_n659), .B2(new_n487), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n717), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n710), .B1(new_n716), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n685), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(new_n680), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n247), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n205), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n674), .B2(G330), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n674), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n209), .A2(new_n311), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n733), .A2(new_n734), .B1(G116), .B2(new_n209), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n242), .A2(new_n285), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n209), .A2(new_n294), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n285), .B2(new_n216), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g0539(.A1(KEYINPUT89), .A2(G13), .A3(G33), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT89), .B1(G13), .B2(G33), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n213), .B1(G20), .B2(new_n307), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n730), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n206), .A2(new_n321), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n362), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n311), .B1(new_n753), .B2(new_n328), .C1(new_n755), .C2(new_n295), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n206), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n303), .A3(new_n362), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n756), .B1(KEYINPUT32), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(KEYINPUT32), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT90), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n763), .B1(new_n769), .B2(G87), .ZN(new_n770));
  OAI21_X1  g0570(.A(G20), .B1(new_n751), .B2(G179), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT91), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G97), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n749), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n303), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n757), .A2(new_n303), .A3(G200), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n249), .B1(new_n781), .B2(new_n378), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n778), .A2(G190), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G68), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n762), .A2(new_n770), .A3(new_n777), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n311), .B1(new_n754), .B2(G311), .ZN(new_n786));
  INV_X1    g0586(.A(new_n758), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G329), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n786), .B(new_n788), .C1(new_n789), .C2(new_n781), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G303), .B2(new_n769), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n775), .A2(new_n476), .B1(new_n792), .B2(new_n780), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT92), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n783), .A2(new_n796), .B1(new_n752), .B2(G322), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n793), .A2(new_n794), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n785), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n748), .B1(new_n801), .B2(new_n745), .ZN(new_n802));
  INV_X1    g0602(.A(new_n744), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n674), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n732), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n374), .A2(new_n656), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n386), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n390), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n616), .A2(new_n657), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n712), .A2(new_n715), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n811), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n647), .A2(new_n657), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n710), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n730), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n812), .A2(new_n710), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n730), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n742), .A2(new_n745), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT94), .Z(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n822), .B2(new_n295), .ZN(new_n823));
  INV_X1    g0623(.A(new_n745), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n754), .A2(G159), .B1(new_n752), .B2(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  INV_X1    g0626(.A(new_n783), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n780), .C1(new_n260), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT34), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n775), .A2(new_n328), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n768), .A2(new_n249), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n758), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n781), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G68), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n311), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n830), .A2(new_n831), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n311), .B1(new_n754), .B2(G116), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n476), .B2(new_n753), .C1(new_n768), .C2(new_n378), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n827), .A2(new_n789), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n781), .A2(new_n222), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  INV_X1    g0642(.A(G311), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n780), .A2(new_n842), .B1(new_n758), .B2(new_n843), .ZN(new_n844));
  NOR4_X1   g0644(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n829), .A2(new_n837), .B1(new_n845), .B2(new_n777), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n823), .B1(new_n824), .B2(new_n846), .C1(new_n813), .C2(new_n743), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n818), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  NOR2_X1   g0649(.A1(new_n727), .A2(new_n205), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT95), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n403), .A2(new_n657), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n440), .A2(new_n441), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n450), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n446), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n613), .A2(new_n614), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n404), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n851), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n442), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n613), .A2(new_n614), .A3(new_n450), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n852), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT95), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n707), .A2(new_n708), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT101), .B1(new_n866), .B2(new_n704), .ZN(new_n867));
  AND4_X1   g0667(.A1(KEYINPUT101), .A2(new_n704), .A3(new_n701), .A4(new_n706), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(new_n811), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT98), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n346), .A2(new_n654), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n625), .B2(new_n622), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n320), .A2(new_n322), .A3(new_n654), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n365), .B1(new_n879), .B2(new_n346), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT97), .B1(new_n358), .B2(new_n878), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n358), .A2(new_n878), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n884), .A2(KEYINPUT97), .A3(KEYINPUT37), .A4(new_n365), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n873), .B(new_n874), .C1(new_n877), .C2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT96), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT16), .B1(new_n356), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n337), .A2(KEYINPUT96), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n348), .B1(new_n891), .B2(new_n357), .ZN(new_n892));
  INV_X1    g0692(.A(new_n654), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n892), .B(new_n893), .C1(new_n361), .C2(new_n369), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n878), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n882), .B1(new_n346), .B2(new_n364), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n895), .A2(new_n896), .B1(new_n880), .B2(new_n882), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n875), .B1(new_n361), .B2(new_n369), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n883), .A3(new_n885), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n873), .B1(new_n901), .B2(new_n874), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n872), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n871), .B1(new_n865), .B2(new_n870), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n894), .A2(new_n897), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n874), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n898), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n865), .A2(new_n870), .A3(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n869), .A2(new_n451), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n915), .A2(new_n916), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n918), .A2(new_n686), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n899), .A2(new_n902), .A3(KEYINPUT39), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n910), .B2(new_n898), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT99), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n874), .B1(new_n877), .B2(new_n886), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT98), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(new_n923), .A3(new_n898), .A4(new_n887), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT99), .ZN(new_n929));
  INV_X1    g0729(.A(new_n911), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n923), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n442), .A2(new_n656), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n814), .A2(new_n810), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n859), .B2(new_n864), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n911), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n361), .A2(new_n654), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n629), .A2(new_n716), .A3(new_n723), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n628), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n850), .B1(new_n921), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n921), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n501), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(G116), .A3(new_n214), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n215), .A2(new_n295), .A3(new_n329), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n220), .A2(G50), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n247), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT103), .ZN(G367));
  OAI21_X1  g0755(.A(new_n746), .B1(new_n209), .B2(new_n573), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n238), .A2(new_n737), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n730), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G143), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n780), .B1(new_n827), .B2(new_n759), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n295), .A2(new_n781), .B1(new_n758), .B2(new_n826), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n311), .B1(new_n753), .B2(new_n260), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G50), .B2(new_n754), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n776), .A2(G68), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n769), .A2(G58), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n294), .B1(new_n753), .B2(new_n842), .C1(new_n755), .C2(new_n789), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n787), .A2(G317), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n780), .B2(new_n843), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n827), .A2(new_n476), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n781), .A2(new_n493), .ZN(new_n972));
  OR4_X1    g0772(.A1(new_n968), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n768), .B2(new_n547), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n378), .C2(new_n775), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n967), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n958), .B1(new_n979), .B2(new_n745), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n595), .A2(new_n656), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n638), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n638), .A2(new_n640), .A3(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n984), .B2(new_n803), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n532), .B1(new_n504), .B2(new_n657), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n531), .A2(new_n528), .A3(new_n656), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n666), .A2(new_n668), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT105), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT105), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n666), .A2(new_n991), .A3(new_n668), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n670), .B2(new_n988), .ZN(new_n997));
  INV_X1    g0797(.A(new_n988), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n669), .A2(KEYINPUT44), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n676), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n995), .A2(new_n1000), .A3(new_n677), .A4(new_n1001), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(KEYINPUT106), .B2(new_n1002), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(KEYINPUT106), .A3(new_n677), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n650), .A2(new_n657), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n671), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(new_n666), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT107), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n675), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n675), .A2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n724), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n724), .B1(new_n1005), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n680), .B(KEYINPUT41), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n729), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n676), .A2(new_n988), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n984), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT43), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n666), .A2(new_n998), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT104), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n986), .A2(new_n488), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n656), .B1(new_n1030), .B2(new_n645), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(KEYINPUT42), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1023), .B(new_n1026), .C1(new_n1029), .C2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1025), .A3(new_n1024), .A4(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1022), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1026), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1023), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1022), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1034), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n985), .B1(new_n1021), .B2(new_n1042), .ZN(G387));
  INV_X1    g0843(.A(new_n1016), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n726), .A3(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n664), .A2(new_n665), .A3(new_n803), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n733), .A2(new_n682), .B1(G107), .B2(new_n209), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n737), .B1(new_n235), .B2(G45), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n285), .B1(new_n220), .B2(new_n295), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT108), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n681), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n265), .A2(KEYINPUT50), .A3(new_n249), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT50), .B1(new_n265), .B2(new_n249), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1052), .B1(new_n1051), .B2(new_n681), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1048), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G283), .A2(new_n776), .B1(new_n769), .B2(G294), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n754), .A2(G303), .B1(new_n752), .B2(G317), .ZN(new_n1058));
  INV_X1    g0858(.A(G322), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n843), .B2(new_n827), .C1(new_n1059), .C2(new_n780), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT110), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT49), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n294), .B1(new_n758), .B2(new_n792), .C1(new_n547), .C2(new_n781), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1066), .B2(KEYINPUT49), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G68), .A2(new_n754), .B1(new_n783), .B2(new_n265), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT109), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n776), .A2(new_n372), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n769), .A2(G77), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n294), .B(new_n972), .C1(G50), .C2(new_n752), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n779), .A2(G159), .B1(new_n787), .B2(G150), .ZN(new_n1075));
  AND4_X1   g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1067), .A2(new_n1069), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n730), .B1(new_n747), .B2(new_n1056), .C1(new_n1077), .C2(new_n824), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1046), .B1(new_n728), .B2(new_n1014), .C1(new_n1047), .C2(new_n1078), .ZN(G393));
  AND2_X1   g0879(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n729), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n998), .A2(new_n744), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT111), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n746), .B1(new_n493), .B2(new_n209), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n245), .A2(new_n737), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n730), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n827), .A2(new_n842), .B1(new_n758), .B2(new_n1059), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n294), .B1(new_n755), .B2(new_n476), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G107), .C2(new_n834), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n779), .B1(new_n752), .B2(G311), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  NAND2_X1  g0891(.A1(new_n776), .A2(G116), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n769), .A2(G283), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n311), .B1(new_n755), .B2(new_n264), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n841), .B(new_n1095), .C1(G50), .C2(new_n783), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G150), .A2(new_n779), .B1(new_n752), .B2(G159), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(new_n295), .C2(new_n775), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n768), .A2(new_n220), .B1(new_n959), .B2(new_n758), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT112), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1094), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1086), .B1(new_n1102), .B2(new_n745), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n726), .B1(new_n1080), .B2(new_n1016), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1005), .A2(new_n1017), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1081), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n932), .B1(new_n934), .B2(new_n938), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n722), .A2(new_n657), .A3(new_n809), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1109), .A2(new_n810), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n859), .B2(new_n864), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT113), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n903), .A2(new_n934), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1109), .A2(new_n810), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT95), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT95), .B1(new_n861), .B2(new_n863), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT113), .B1(new_n1119), .B2(new_n1113), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1108), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(G330), .B(new_n813), .C1(new_n867), .C2(new_n868), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n859), .B2(new_n864), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(KEYINPUT114), .A3(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n686), .B(new_n811), .C1(new_n705), .C2(new_n709), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n865), .B(new_n1125), .C1(KEYINPUT114), .C2(new_n1122), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1108), .B(new_n1126), .C1(new_n1115), .C2(new_n1120), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n729), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n819), .B1(new_n822), .B2(new_n264), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n780), .A2(new_n789), .B1(new_n758), .B2(new_n476), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n835), .B1(new_n753), .B2(new_n547), .C1(new_n755), .C2(new_n493), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1130), .B(new_n1131), .C1(G107), .C2(new_n783), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n294), .B1(new_n768), .B2(new_n222), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT118), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(new_n295), .C2(new_n775), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n768), .A2(new_n260), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n311), .B1(new_n753), .B2(new_n832), .C1(new_n755), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1140), .A2(new_n780), .B1(new_n827), .B2(new_n826), .ZN(new_n1141));
  INV_X1    g0941(.A(G125), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n249), .A2(new_n781), .B1(new_n758), .B2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1137), .B(new_n1144), .C1(new_n759), .C2(new_n775), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1135), .A2(new_n1145), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1129), .B1(new_n824), .B2(new_n1146), .C1(new_n933), .C2(new_n743), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1112), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1119), .A2(KEYINPUT113), .A3(new_n1113), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n934), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n937), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1149), .A2(new_n1150), .B1(new_n1153), .B2(new_n932), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1123), .A2(KEYINPUT114), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1127), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1116), .B1(new_n865), .B2(new_n1125), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT115), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1122), .A2(new_n859), .A3(new_n1158), .A4(new_n864), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1122), .A2(new_n859), .A3(new_n864), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT115), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1157), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n865), .A2(new_n1125), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n936), .B1(new_n1163), .B2(new_n1123), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n629), .B(G330), .C1(new_n867), .C2(new_n868), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n627), .A2(new_n1166), .A3(new_n309), .A4(new_n942), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1148), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1124), .A2(KEYINPUT116), .A3(new_n1127), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n680), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1156), .A2(new_n1169), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1173), .A2(KEYINPUT117), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1128), .B(new_n1147), .C1(new_n1176), .C2(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n268), .A2(new_n893), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n310), .B(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1181), .B(new_n1182), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n908), .A2(G330), .A3(new_n914), .A4(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n914), .B(G330), .C1(new_n906), .C2(new_n907), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1183), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n941), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n941), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1185), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1167), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(KEYINPUT119), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT119), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1195), .B(new_n1167), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1179), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1168), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1195), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(KEYINPUT119), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(KEYINPUT57), .A3(new_n1192), .A4(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1202), .A3(new_n726), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1183), .A2(new_n742), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n742), .A2(G50), .A3(new_n745), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n311), .A2(new_n480), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G50), .B(new_n1206), .C1(new_n262), .C2(new_n281), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n780), .A2(new_n547), .B1(new_n781), .B2(new_n328), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n827), .A2(new_n493), .B1(new_n758), .B2(new_n789), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1206), .B1(new_n753), .B2(new_n378), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n372), .B2(new_n754), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1212), .A3(new_n965), .A4(new_n1073), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n754), .A2(G137), .B1(new_n752), .B2(G128), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1142), .B2(new_n780), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G132), .B2(new_n783), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n260), .B2(new_n775), .C1(new_n768), .C2(new_n1138), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n262), .B(new_n281), .C1(new_n781), .C2(new_n759), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G124), .B2(new_n787), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1215), .B1(new_n1214), .B2(new_n1213), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n819), .B(new_n1205), .C1(new_n1225), .C2(new_n745), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1192), .A2(new_n729), .B1(new_n1204), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1203), .A2(new_n1227), .ZN(G375));
  NAND3_X1  g1028(.A1(new_n1162), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1169), .A2(new_n1020), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n819), .B1(new_n822), .B2(new_n220), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n294), .B1(new_n754), .B2(G150), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n826), .B2(new_n753), .C1(new_n768), .C2(new_n759), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n775), .A2(new_n249), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n827), .A2(new_n1138), .B1(new_n328), .B2(new_n781), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n780), .A2(new_n832), .B1(new_n758), .B2(new_n1140), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1072), .B1(new_n789), .B2(new_n753), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT120), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n779), .A2(G294), .B1(new_n787), .B2(G303), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n547), .B2(new_n827), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n294), .B1(new_n295), .B2(new_n781), .C1(new_n755), .C2(new_n378), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G97), .C2(new_n769), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1237), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1231), .B1(new_n824), .B2(new_n1244), .C1(new_n865), .C2(new_n743), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1165), .B2(new_n729), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1230), .A2(new_n1247), .ZN(G381));
  OR4_X1    g1048(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(G387), .A3(G381), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1128), .A2(new_n1147), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1177), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1254), .A3(new_n1227), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1055(.A1(new_n655), .A2(G213), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(G375), .A2(G378), .A3(new_n1256), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT121), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G213), .A3(G407), .ZN(G409));
  NAND3_X1  g1059(.A1(new_n1203), .A2(G378), .A3(new_n1227), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1227), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1194), .A2(new_n1196), .A3(new_n1019), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1254), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1256), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1229), .B1(new_n1171), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1162), .A2(new_n1164), .A3(KEYINPUT60), .A4(new_n1167), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n726), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT122), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1267), .A2(KEYINPUT122), .A3(new_n726), .A4(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1247), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n848), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(G384), .A3(new_n1247), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(KEYINPUT123), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1273), .B2(new_n1247), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1247), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n848), .B(new_n1280), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1278), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n655), .A2(G213), .A3(G2897), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1284), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1286), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1265), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1264), .A2(new_n1256), .A3(new_n1283), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT62), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1264), .A2(new_n1297), .A3(new_n1256), .A4(new_n1283), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1293), .A2(new_n1295), .A3(new_n1296), .A4(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n805), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G390), .B(new_n985), .C1(new_n1021), .C2(new_n1042), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1301), .B1(new_n1305), .B2(KEYINPUT125), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1307), .B(new_n1300), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1299), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1309), .B2(new_n1296), .ZN(new_n1313));
  NOR4_X1   g1113(.A1(new_n1306), .A2(new_n1308), .A3(KEYINPUT126), .A4(KEYINPUT61), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1294), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1294), .A2(new_n1316), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1315), .A2(new_n1317), .A3(new_n1293), .A4(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1319), .ZN(G405));
  OR2_X1    g1120(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1254), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1322), .B(new_n1260), .C1(new_n1279), .C2(new_n1281), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1260), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1283), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1321), .A2(new_n1323), .A3(new_n1325), .A4(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1325), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1323), .ZN(new_n1329));
  OAI211_X1 g1129(.A(KEYINPUT127), .B(new_n1310), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(G402));
endmodule


