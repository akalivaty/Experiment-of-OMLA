//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1182, new_n1183,
    new_n1184, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G238), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n203), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n206), .B1(KEYINPUT1), .B2(new_n215), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XOR2_X1   g0023(.A(G238), .B(G244), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n225), .B(new_n226), .Z(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XOR2_X1   g0031(.A(G68), .B(G77), .Z(new_n232));
  XOR2_X1   g0032(.A(G50), .B(G58), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G351));
  OR2_X1    g0038(.A1(KEYINPUT66), .A2(G1), .ZN(new_n239));
  NAND2_X1  g0039(.A1(KEYINPUT66), .A2(G1), .ZN(new_n240));
  NAND4_X1  g0040(.A1(new_n239), .A2(G13), .A3(G20), .A4(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT69), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g0043(.A1(KEYINPUT66), .A2(G1), .ZN(new_n244));
  NOR2_X1   g0044(.A1(KEYINPUT66), .A2(G1), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n246), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n216), .B1(new_n203), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n246), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G50), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n243), .A2(new_n247), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n258), .A3(new_n208), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n259), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT68), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n256), .A2(new_n257), .B1(new_n266), .B2(new_n250), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n255), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n239), .A2(new_n240), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G41), .A2(G45), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT67), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G226), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n217), .B2(new_n269), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1698), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(G222), .B2(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n275), .B(new_n279), .C1(new_n270), .C2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n268), .A2(KEYINPUT9), .B1(new_n291), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n292), .B1(KEYINPUT9), .B2(new_n268), .C1(new_n293), .C2(new_n291), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n268), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G179), .B2(new_n291), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n257), .A2(new_n208), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n264), .B2(new_n283), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n250), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT11), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G97), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n249), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n289), .B2(G226), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n270), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n312), .A2(new_n313), .B1(new_n277), .B2(new_n278), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n274), .A2(G238), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(G169), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n321), .B1(new_n320), .B2(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n307), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n307), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n317), .A2(G190), .A3(new_n319), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n320), .A2(G200), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT70), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AND4_X1   g0131(.A1(KEYINPUT70), .A2(new_n330), .A3(new_n328), .A4(new_n327), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n265), .A2(G20), .A3(G33), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n336), .A2(new_n263), .B1(new_n262), .B2(new_n283), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n250), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n334), .B(new_n338), .C1(G77), .C2(new_n248), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n289), .A2(G232), .B1(G107), .B2(new_n288), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n207), .B2(new_n281), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n313), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n274), .A2(G244), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n279), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n339), .B1(G200), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n293), .B2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n296), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n339), .C1(G179), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n299), .A2(new_n333), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n265), .B1(G20), .B2(new_n246), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT74), .ZN(new_n352));
  INV_X1    g0152(.A(new_n265), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n352), .A2(new_n252), .B1(new_n248), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n258), .A2(new_n208), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n286), .A2(KEYINPUT72), .A3(G33), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n285), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT72), .B1(new_n286), .B2(G33), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT7), .B(new_n262), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G20), .B2(new_n280), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n208), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT73), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n359), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT73), .B(new_n208), .C1(new_n363), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n355), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n262), .A3(new_n288), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT7), .B1(new_n280), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G68), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n359), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n250), .B1(new_n374), .B2(new_n355), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n354), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(G232), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n279), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n285), .A2(new_n287), .A3(G226), .A4(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n280), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  INV_X1    g0184(.A(G1698), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n280), .A2(G223), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n379), .B1(new_n387), .B2(new_n313), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G179), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n296), .B2(new_n388), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n377), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT18), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  AOI211_X1 g0194(.A(G190), .B(new_n379), .C1(new_n313), .C2(new_n387), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n387), .A2(new_n313), .ZN(new_n396));
  INV_X1    g0196(.A(new_n379), .ZN(new_n397));
  AOI21_X1  g0197(.A(G200), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n397), .A3(new_n293), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(KEYINPUT76), .C1(G200), .C2(new_n388), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n377), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT77), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT77), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n405), .A3(new_n377), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n404), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n402), .A2(new_n405), .A3(new_n377), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n402), .B2(new_n377), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n403), .B2(KEYINPUT17), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n393), .B(new_n407), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n350), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G283), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n262), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT79), .B(G97), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n249), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT20), .ZN(new_n422));
  INV_X1    g0222(.A(G116), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G20), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n250), .A2(new_n424), .ZN(new_n425));
  OR3_X1    g0225(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n422), .B1(new_n421), .B2(new_n425), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n257), .B2(new_n423), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n246), .A2(G33), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n248), .A2(G116), .A3(new_n251), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT5), .B(G41), .Z(new_n433));
  NAND3_X1  g0233(.A1(new_n239), .A2(G45), .A3(new_n240), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n313), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(G270), .B1(new_n277), .B2(new_n435), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n280), .A2(G264), .A3(G1698), .ZN(new_n438));
  INV_X1    g0238(.A(G303), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n280), .A2(G257), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n438), .B1(new_n439), .B2(new_n280), .C1(new_n440), .C2(G1698), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n313), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n432), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n431), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n431), .B2(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n437), .A2(new_n442), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n293), .C2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n296), .B1(new_n437), .B2(new_n442), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n431), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT21), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n431), .A2(new_n449), .A3(KEYINPUT21), .ZN(new_n453));
  INV_X1    g0253(.A(G179), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n431), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n280), .A2(G250), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n280), .A2(KEYINPUT83), .A3(G250), .A4(new_n385), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G294), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n440), .A2(new_n385), .B1(new_n249), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n270), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n435), .A2(new_n277), .ZN(new_n469));
  OAI211_X1 g0269(.A(G264), .B(new_n270), .C1(new_n433), .C2(new_n434), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G190), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n280), .A2(new_n262), .A3(G87), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT22), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G20), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT23), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G116), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n478), .A2(KEYINPUT23), .B1(G20), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n478), .B2(KEYINPUT23), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n475), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n476), .B1(new_n475), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n250), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n248), .A2(new_n251), .A3(new_n429), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n257), .A2(KEYINPUT25), .A3(new_n477), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT25), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n248), .B2(G107), .ZN(new_n492));
  AOI22_X1  g0292(.A1(G107), .A2(new_n489), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n471), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n466), .B1(new_n462), .B2(new_n463), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(new_n270), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n473), .A2(new_n488), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n308), .A2(new_n477), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g0301(.A(KEYINPUT79), .B(G97), .Z(new_n502));
  NAND2_X1  g0302(.A1(new_n477), .A2(KEYINPUT6), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n501), .A2(KEYINPUT6), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n363), .A2(new_n365), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G107), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n250), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n248), .A2(G97), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n489), .B2(G97), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n288), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n385), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n418), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n385), .B1(new_n461), .B2(KEYINPUT4), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n313), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n436), .A2(G257), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n469), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n509), .A2(new_n511), .B1(new_n520), .B2(new_n296), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n454), .A3(new_n469), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(G190), .A3(new_n469), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(G200), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n509), .A3(new_n511), .A4(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n498), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n488), .A2(new_n493), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n296), .B1(new_n468), .B2(new_n471), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n494), .B(new_n454), .C1(new_n495), .C2(new_n270), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n502), .B2(new_n263), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n280), .A2(new_n262), .A3(G68), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n420), .A2(G87), .A3(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(new_n309), .B2(KEYINPUT19), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n250), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n257), .A2(new_n336), .ZN(new_n540));
  INV_X1    g0340(.A(new_n336), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n248), .A2(new_n251), .A3(new_n541), .A4(new_n429), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n280), .A2(G244), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n280), .A2(G238), .A3(new_n385), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n482), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n313), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n270), .A2(G274), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT80), .B1(new_n548), .B2(new_n434), .ZN(new_n549));
  INV_X1    g0349(.A(G45), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n244), .A2(new_n245), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT80), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n277), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n434), .A2(G250), .A3(new_n270), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n547), .A2(new_n554), .A3(new_n454), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n547), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n555), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n543), .B(new_n556), .C1(new_n559), .C2(G169), .ZN(new_n560));
  OAI21_X1  g0360(.A(G200), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n538), .A2(new_n250), .B1(new_n257), .B2(new_n336), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n489), .A2(G87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n547), .A2(new_n554), .A3(G190), .A4(new_n555), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n532), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AND4_X1   g0366(.A1(new_n417), .A2(new_n459), .A3(new_n528), .A4(new_n566), .ZN(G372));
  NOR2_X1   g0367(.A1(new_n331), .A2(new_n332), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n348), .A2(KEYINPUT87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n348), .A2(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n326), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n407), .C1(new_n411), .C2(new_n413), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n393), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n295), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(new_n298), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n563), .A2(new_n562), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n559), .B2(G190), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n554), .A2(KEYINPUT84), .A3(new_n555), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n557), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT85), .B1(new_n582), .B2(new_n432), .ZN(new_n583));
  INV_X1    g0383(.A(new_n581), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT84), .B1(new_n554), .B2(new_n555), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n547), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(G200), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n578), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n556), .B(new_n543), .C1(new_n582), .C2(G169), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT26), .ZN(new_n592));
  INV_X1    g0392(.A(new_n524), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n590), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n521), .A2(new_n560), .A3(new_n523), .A4(new_n565), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(KEYINPUT26), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(KEYINPUT86), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n530), .A2(new_n531), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n488), .B2(new_n493), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n591), .B(new_n528), .C1(new_n457), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT86), .B1(new_n594), .B2(new_n597), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n417), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n576), .A2(new_n605), .ZN(G369));
  INV_X1    g0406(.A(G13), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n246), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G213), .B1(new_n609), .B2(KEYINPUT27), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(KEYINPUT27), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G343), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n431), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n459), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n458), .B2(new_n619), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G330), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n529), .A2(new_n618), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n600), .B1(new_n624), .B2(new_n498), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n532), .A2(new_n618), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n626), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n458), .A2(new_n618), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(G399));
  NAND2_X1  g0432(.A1(new_n536), .A2(new_n423), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n204), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G41), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(G1), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n219), .B2(new_n637), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT28), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n457), .B2(new_n600), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n450), .A2(new_n451), .B1(new_n455), .B2(new_n431), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n532), .A2(new_n643), .A3(KEYINPUT90), .A4(new_n453), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n591), .A2(new_n642), .A3(new_n528), .A4(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n590), .B1(new_n596), .B2(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n593), .A2(new_n589), .A3(new_n590), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(KEYINPUT26), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(KEYINPUT89), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n650), .B(new_n646), .C1(KEYINPUT26), .C2(new_n647), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT29), .B1(new_n652), .B2(new_n618), .ZN(new_n653));
  INV_X1    g0453(.A(new_n618), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n604), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(KEYINPUT29), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n522), .A2(new_n559), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n455), .A3(new_n472), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT30), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(G179), .B1(new_n437), .B2(new_n442), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n586), .A2(new_n520), .A3(new_n496), .A4(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n658), .A2(KEYINPUT30), .A3(new_n455), .A4(new_n472), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n618), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT31), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(KEYINPUT31), .A3(new_n618), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n459), .A2(new_n528), .A3(new_n566), .A4(new_n654), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n657), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n640), .B1(new_n673), .B2(G1), .ZN(G364));
  INV_X1    g0474(.A(G1), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n608), .B2(G45), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n637), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n623), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(G330), .B2(new_n621), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n280), .A2(new_n204), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(KEYINPUT91), .B2(G355), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(KEYINPUT91), .B2(G355), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(G116), .B2(new_n204), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n234), .A2(G45), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n635), .A2(new_n280), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n220), .B2(new_n550), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G13), .A2(G33), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G20), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n216), .B1(G20), .B2(new_n296), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n678), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n262), .A2(new_n293), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n454), .A3(G200), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT94), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n454), .A2(G200), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n262), .A2(G190), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n702), .A2(G87), .B1(G77), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n704), .A2(new_n454), .A3(new_n432), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G159), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n697), .A2(new_n703), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  OAI221_X1 g0515(.A(new_n710), .B1(KEYINPUT32), .B2(new_n713), .C1(new_n258), .C2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n262), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n308), .ZN(new_n719));
  NAND3_X1  g0519(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G190), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(G68), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n720), .A2(new_n293), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G50), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n713), .A2(KEYINPUT32), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n704), .A2(new_n454), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n477), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n288), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n722), .A2(new_n724), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n714), .ZN(new_n730));
  XNOR2_X1  g0530(.A(KEYINPUT33), .B(G317), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n730), .A2(G322), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NAND2_X1  g0533(.A1(new_n702), .A2(G303), .ZN(new_n734));
  INV_X1    g0534(.A(new_n723), .ZN(new_n735));
  INV_X1    g0535(.A(G326), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n718), .A2(new_n465), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(G329), .B2(new_n712), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n709), .A2(G311), .ZN(new_n739));
  INV_X1    g0539(.A(new_n726), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n280), .B1(new_n740), .B2(G283), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n716), .A2(new_n729), .B1(new_n733), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n696), .B1(new_n743), .B2(new_n693), .ZN(new_n744));
  INV_X1    g0544(.A(new_n692), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n621), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n680), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(G396));
  NAND4_X1  g0548(.A1(new_n569), .A2(new_n339), .A3(new_n570), .A4(new_n618), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n618), .A2(new_n339), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n346), .A2(new_n348), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n655), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n654), .B(new_n752), .C1(new_n602), .C2(new_n603), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n672), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n637), .B2(new_n676), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n672), .A3(new_n755), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n693), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n721), .A2(G150), .B1(new_n723), .B2(G137), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  INV_X1    g0562(.A(G143), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n761), .B1(new_n708), .B2(new_n762), .C1(new_n715), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT34), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n280), .B1(new_n726), .B2(new_n208), .ZN(new_n766));
  INV_X1    g0566(.A(G132), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n718), .A2(new_n258), .B1(new_n711), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n766), .B(new_n768), .C1(new_n702), .C2(G50), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G87), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n726), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n721), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n773), .A2(new_n774), .B1(new_n735), .B2(new_n439), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(G311), .C2(new_n712), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n702), .A2(G107), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n709), .A2(G116), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n280), .B(new_n719), .C1(G294), .C2(new_n730), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n760), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n693), .A2(new_n690), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n677), .B(new_n781), .C1(new_n283), .C2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n752), .B2(new_n691), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n759), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G384));
  OAI21_X1  g0586(.A(G77), .B1(new_n258), .B2(new_n208), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n787), .A2(new_n219), .B1(G50), .B2(new_n208), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n607), .A3(new_n271), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n423), .B(new_n218), .C1(new_n504), .C2(KEYINPUT35), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(KEYINPUT35), .B2(new_n504), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT36), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT40), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n375), .B1(new_n355), .B2(new_n374), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(new_n354), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(new_n615), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n414), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n390), .B2(new_n615), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n404), .A2(new_n801), .A3(new_n406), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT37), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n408), .A2(new_n409), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n377), .A2(new_n616), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n392), .A2(new_n805), .A3(KEYINPUT37), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n800), .A2(KEYINPUT38), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(KEYINPUT97), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT97), .ZN(new_n814));
  AOI221_X4 g0614(.A(new_n810), .B1(new_n803), .B2(new_n807), .C1(new_n414), .C2(new_n799), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT38), .B1(new_n800), .B2(new_n808), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n307), .A2(new_n618), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n333), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n326), .B(new_n819), .C1(new_n331), .C2(new_n332), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n753), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n670), .A2(KEYINPUT101), .A3(new_n671), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n671), .A2(new_n669), .A3(new_n668), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT101), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n823), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n796), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT102), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n370), .A2(new_n376), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n390), .B1(new_n832), .B2(new_n354), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n615), .B1(new_n832), .B2(new_n354), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(new_n403), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(KEYINPUT98), .B1(new_n804), .B2(new_n806), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n414), .A2(new_n805), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT38), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n831), .B1(new_n841), .B2(new_n815), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n837), .A2(new_n838), .B1(new_n414), .B2(new_n805), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n812), .B(KEYINPUT102), .C1(new_n843), .C2(KEYINPUT38), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n830), .A2(new_n842), .A3(KEYINPUT40), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n829), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n824), .A2(new_n827), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n416), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n846), .A2(new_n848), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n850), .A2(new_n657), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n326), .A2(new_n618), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT39), .B1(new_n815), .B2(new_n816), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n812), .B(new_n855), .C1(new_n843), .C2(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT100), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(KEYINPUT100), .A3(new_n856), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n853), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n821), .A2(new_n822), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n348), .A2(new_n618), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n863), .B1(new_n755), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n818), .A2(new_n867), .B1(new_n393), .B2(new_n615), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n656), .A2(new_n417), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n871), .A2(new_n576), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n852), .A2(new_n873), .B1(new_n246), .B2(new_n608), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n852), .A2(new_n873), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n795), .B1(new_n874), .B2(new_n875), .ZN(G367));
  OAI221_X1 g0676(.A(new_n694), .B1(new_n204), .B2(new_n336), .C1(new_n230), .C2(new_n687), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(new_n678), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n618), .A2(new_n577), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n590), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT103), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n591), .A2(new_n879), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT104), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n701), .A2(new_n423), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT46), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n708), .A2(new_n774), .B1(new_n477), .B2(new_n718), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT108), .Z(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT109), .B(G311), .Z(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n723), .B1(G294), .B2(new_n721), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n502), .B2(new_n726), .ZN(new_n891));
  INV_X1    g0691(.A(G317), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n288), .B1(new_n892), .B2(new_n711), .C1(new_n715), .C2(new_n439), .ZN(new_n893));
  NOR4_X1   g0693(.A1(new_n886), .A2(new_n888), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT110), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT110), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n726), .A2(new_n283), .ZN(new_n898));
  INV_X1    g0698(.A(G150), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n280), .B1(new_n714), .B2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n898), .B(new_n900), .C1(new_n702), .C2(G58), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n718), .A2(new_n208), .ZN(new_n902));
  INV_X1    g0702(.A(G137), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n773), .A2(new_n762), .B1(new_n711), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n902), .B(new_n904), .C1(G143), .C2(new_n723), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n901), .B(new_n905), .C1(new_n256), .C2(new_n708), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT111), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n896), .A2(new_n897), .A3(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT47), .Z(new_n909));
  OAI221_X1 g0709(.A(new_n878), .B1(new_n884), .B2(new_n745), .C1(new_n760), .C2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n593), .A2(new_n618), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n509), .A2(new_n511), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n524), .B(new_n527), .C1(new_n913), .C2(new_n654), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n631), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n524), .B1(new_n914), .B2(new_n532), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n654), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n911), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT105), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(new_n911), .C2(new_n921), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n628), .A2(new_n916), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n927), .B(new_n928), .Z(new_n929));
  XNOR2_X1  g0729(.A(new_n676), .B(KEYINPUT107), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n631), .A2(new_n629), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n916), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT44), .Z(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n916), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT45), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n628), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n627), .B(new_n630), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n622), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n628), .A3(new_n936), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n673), .A2(new_n939), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n673), .ZN(new_n945));
  XOR2_X1   g0745(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n946));
  XNOR2_X1  g0746(.A(new_n636), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n931), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n910), .B1(new_n929), .B2(new_n949), .ZN(G387));
  OAI21_X1  g0750(.A(new_n941), .B1(new_n656), .B2(new_n672), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n673), .A2(new_n942), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n952), .A2(new_n636), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(G45), .B(new_n633), .C1(G68), .C2(G77), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT113), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n265), .A2(KEYINPUT50), .A3(G50), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT50), .B1(new_n265), .B2(G50), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n957), .A2(KEYINPUT113), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n686), .B1(new_n550), .B2(new_n227), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n634), .A2(new_n681), .B1(G107), .B2(new_n204), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT112), .Z(new_n965));
  AND2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n678), .B1(new_n966), .B2(new_n695), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n889), .A2(new_n721), .B1(G322), .B2(new_n723), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n708), .B2(new_n439), .C1(new_n715), .C2(new_n892), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT48), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  INV_X1    g0772(.A(new_n718), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n702), .A2(G294), .B1(G283), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(KEYINPUT49), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n288), .B1(new_n711), .B2(new_n736), .C1(new_n423), .C2(new_n726), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(KEYINPUT49), .B2(new_n976), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n718), .A2(new_n336), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n735), .A2(new_n762), .B1(new_n726), .B2(new_n308), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n353), .C2(new_n721), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n280), .B1(new_n714), .B2(new_n256), .C1(new_n899), .C2(new_n711), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n709), .B2(G68), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(new_n283), .C2(new_n701), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n967), .B1(new_n987), .B2(new_n693), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n627), .A2(new_n745), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n942), .B2(new_n931), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n955), .A2(new_n994), .ZN(G393));
  OR2_X1    g0795(.A1(new_n943), .A2(KEYINPUT116), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n943), .A2(KEYINPUT116), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n939), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n953), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n636), .A3(new_n944), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n694), .B1(new_n204), .B2(new_n502), .C1(new_n237), .C2(new_n687), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n678), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n288), .B(new_n772), .C1(new_n709), .C2(new_n353), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n735), .A2(new_n899), .B1(new_n714), .B2(new_n762), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT51), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n702), .A2(G68), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n773), .A2(new_n256), .B1(new_n711), .B2(new_n763), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G77), .B2(new_n973), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n280), .B(new_n727), .C1(new_n709), .C2(G294), .ZN(new_n1010));
  INV_X1    g0810(.A(G322), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n773), .A2(new_n439), .B1(new_n711), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G116), .B2(new_n973), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1010), .B(new_n1013), .C1(new_n774), .C2(new_n701), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n730), .A2(G311), .B1(new_n723), .B2(G317), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT52), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1009), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1002), .B1(new_n1017), .B2(new_n693), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n915), .B2(new_n745), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1000), .B(new_n1019), .C1(new_n930), .C2(new_n998), .ZN(G390));
  NAND3_X1  g0820(.A1(new_n824), .A2(new_n827), .A3(G330), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n823), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n867), .A2(new_n853), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n859), .A2(new_n860), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n853), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n654), .B(new_n752), .C1(new_n649), .C2(new_n651), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n865), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n821), .A2(new_n822), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n842), .A3(new_n844), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1023), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT117), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n854), .A2(KEYINPUT100), .A3(new_n856), .ZN(new_n1034));
  AOI21_X1  g0834(.A(KEYINPUT100), .B1(new_n854), .B2(new_n856), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n866), .A2(new_n1026), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n672), .A2(new_n752), .A3(new_n1029), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1033), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1041), .A2(new_n1025), .A3(KEYINPUT117), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1032), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n672), .A2(new_n752), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1023), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n755), .A2(new_n865), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n863), .B1(new_n1021), .B2(new_n753), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1028), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1045), .A2(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n416), .A2(new_n1021), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n871), .A2(new_n576), .A3(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n636), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1023), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g0856(.A1(new_n1037), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT117), .B1(new_n1041), .B2(new_n1025), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1052), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT118), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1052), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT118), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n636), .A4(new_n1059), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1034), .A2(new_n1035), .A3(new_n691), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n677), .B1(new_n265), .B2(new_n782), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n721), .A2(G107), .B1(new_n723), .B2(G283), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n283), .B2(new_n718), .C1(new_n465), .C2(new_n711), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n280), .B1(new_n730), .B2(G116), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n208), .B2(new_n726), .C1(new_n701), .C2(new_n771), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n420), .C2(new_n709), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n701), .A2(new_n899), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n280), .B1(new_n726), .B2(new_n256), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT119), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n712), .A2(G125), .B1(new_n730), .B2(G132), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT54), .B(G143), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n708), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(G128), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n735), .A2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n718), .A2(new_n762), .B1(new_n773), .B2(new_n903), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1074), .B1(new_n1077), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1069), .B1(new_n1087), .B2(new_n760), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1062), .A2(new_n930), .B1(new_n1068), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1067), .A2(new_n1090), .ZN(G378));
  INV_X1    g0891(.A(G41), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n288), .C1(new_n714), .C2(new_n477), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n902), .B(new_n1093), .C1(new_n702), .C2(G77), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n726), .A2(new_n258), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n773), .A2(new_n308), .B1(new_n735), .B2(new_n423), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G283), .C2(new_n712), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1094), .B(new_n1097), .C1(new_n336), .C2(new_n708), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT58), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(G50), .B1(new_n249), .B2(new_n1092), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n280), .B2(G41), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n773), .A2(new_n767), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n718), .A2(new_n899), .B1(new_n714), .B2(new_n1083), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G125), .C2(new_n723), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n903), .B2(new_n708), .C1(new_n701), .C2(new_n1081), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT59), .Z(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n740), .A2(G159), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G33), .B(G41), .C1(new_n712), .C2(G124), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1108), .A2(KEYINPUT121), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1103), .B1(new_n1099), .B2(new_n1098), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n693), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT122), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n677), .B1(new_n256), .B2(new_n782), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT123), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n268), .A2(new_n616), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT124), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n299), .B(new_n1121), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1123));
  XNOR2_X1  g0923(.A(new_n1122), .B(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1116), .B(new_n1119), .C1(new_n1124), .C2(new_n690), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n861), .A2(new_n868), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n829), .A2(G330), .A3(new_n845), .A4(new_n1124), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n828), .B1(new_n813), .B2(new_n817), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n845), .B(G330), .C1(new_n1128), .C2(KEYINPUT40), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1124), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1127), .A2(new_n1131), .B1(new_n862), .B2(new_n869), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1125), .B1(new_n1134), .B2(new_n931), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1051), .B(KEYINPUT125), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n870), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(KEYINPUT57), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n636), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1136), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1059), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT57), .B1(new_n1144), .B2(new_n1134), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1135), .B1(new_n1142), .B2(new_n1145), .ZN(G375));
  OAI22_X1  g0946(.A1(new_n773), .A2(new_n423), .B1(new_n735), .B2(new_n465), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n981), .B(new_n1147), .C1(G303), .C2(new_n712), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n709), .A2(G107), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n702), .A2(G97), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n280), .B(new_n898), .C1(G283), .C2(new_n730), .ZN(new_n1151));
  AND4_X1   g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n701), .A2(new_n762), .B1(new_n715), .B2(new_n903), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n280), .B1(new_n258), .B2(new_n726), .C1(new_n708), .C2(new_n899), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n718), .A2(new_n256), .B1(new_n735), .B2(new_n767), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n773), .A2(new_n1081), .B1(new_n711), .B2(new_n1083), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n693), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n677), .B1(new_n208), .B2(new_n782), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n1029), .C2(new_n691), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1049), .B2(new_n930), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1063), .A2(new_n948), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1049), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1051), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1162), .B1(new_n1163), .B2(new_n1166), .ZN(G381));
  OR2_X1    g0967(.A1(G387), .A2(G390), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n955), .A2(new_n747), .A3(new_n994), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1168), .A2(G384), .A3(G381), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1125), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n930), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n1132), .A2(new_n1133), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n637), .B1(new_n1175), .B2(new_n1144), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1137), .B2(new_n1172), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n637), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1089), .B1(new_n1059), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1170), .A2(new_n1178), .A3(new_n1180), .ZN(G407));
  NAND2_X1  g0981(.A1(new_n617), .A2(G213), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(G407), .A2(G213), .A3(new_n1184), .ZN(G409));
  NAND3_X1  g0985(.A1(new_n1144), .A2(new_n1134), .A3(new_n948), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1135), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1180), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1089), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(G375), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1164), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT60), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n636), .B(new_n1063), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(G384), .A3(new_n1162), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G384), .B1(new_n1194), .B2(new_n1162), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n1182), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT62), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT61), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT62), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1190), .A2(new_n1202), .A3(new_n1182), .A4(new_n1198), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1197), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n1195), .A3(G2897), .A4(new_n1183), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1183), .A2(G2897), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G378), .A2(new_n1178), .B1(new_n1180), .B2(new_n1187), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n1183), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G387), .A2(G390), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1168), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G393), .A2(G396), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1214), .A2(new_n1169), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1168), .A2(new_n1217), .A3(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1199), .A2(KEYINPUT63), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT63), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1190), .A2(new_n1222), .A3(new_n1182), .A4(new_n1198), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT126), .B1(new_n1209), .B2(new_n1183), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT126), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1190), .A2(new_n1226), .A3(new_n1182), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1227), .A3(new_n1208), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1219), .A2(KEYINPUT61), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1224), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1220), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT127), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1220), .A2(new_n1230), .A3(KEYINPUT127), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(G405));
  NAND2_X1  g1035(.A1(G375), .A2(new_n1180), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1189), .B2(G375), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(new_n1198), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(new_n1219), .ZN(G402));
endmodule


