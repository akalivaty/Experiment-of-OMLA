

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740;

  NAND2_X1 U376 ( .A1(n388), .A2(n386), .ZN(n549) );
  AND2_X2 U377 ( .A1(n391), .A2(n389), .ZN(n388) );
  AND2_X2 U378 ( .A1(n602), .A2(n398), .ZN(n383) );
  INV_X1 U379 ( .A(G953), .ZN(n727) );
  NOR2_X1 U380 ( .A1(n663), .A2(n561), .ZN(n632) );
  NAND2_X1 U381 ( .A1(n393), .A2(n394), .ZN(n507) );
  XNOR2_X1 U382 ( .A(n418), .B(n471), .ZN(n619) );
  XNOR2_X1 U383 ( .A(G146), .B(KEYINPUT4), .ZN(n371) );
  NOR2_X1 U384 ( .A1(n735), .A2(n567), .ZN(n568) );
  XNOR2_X1 U385 ( .A(n558), .B(KEYINPUT105), .ZN(n735) );
  NOR2_X1 U386 ( .A1(n554), .A2(n576), .ZN(n555) );
  XNOR2_X1 U387 ( .A(n413), .B(n412), .ZN(n739) );
  XNOR2_X1 U388 ( .A(n530), .B(n367), .ZN(n734) );
  XOR2_X1 U389 ( .A(n507), .B(KEYINPUT38), .Z(n672) );
  NOR2_X1 U390 ( .A1(n556), .A2(n574), .ZN(n364) );
  NAND2_X1 U391 ( .A1(n399), .A2(n397), .ZN(n396) );
  OR2_X1 U392 ( .A1(n619), .A2(n385), .ZN(n399) );
  INV_X1 U393 ( .A(n477), .ZN(n385) );
  NAND2_X1 U394 ( .A1(n477), .A2(n398), .ZN(n397) );
  NAND2_X1 U395 ( .A1(n671), .A2(KEYINPUT19), .ZN(n392) );
  XNOR2_X1 U396 ( .A(n371), .B(n370), .ZN(n443) );
  AND2_X1 U397 ( .A1(n566), .A2(n565), .ZN(n420) );
  NAND2_X1 U398 ( .A1(n365), .A2(n364), .ZN(n558) );
  XNOR2_X2 U399 ( .A(n363), .B(KEYINPUT22), .ZN(n576) );
  OR2_X1 U400 ( .A1(G902), .A2(G237), .ZN(n478) );
  NAND2_X1 U401 ( .A1(n619), .A2(n395), .ZN(n394) );
  XNOR2_X1 U402 ( .A(n444), .B(G101), .ZN(n445) );
  INV_X1 U403 ( .A(KEYINPUT65), .ZN(n444) );
  XOR2_X1 U404 ( .A(KEYINPUT68), .B(G137), .Z(n460) );
  XOR2_X1 U405 ( .A(n436), .B(KEYINPUT10), .Z(n481) );
  XNOR2_X1 U406 ( .A(G125), .B(G140), .ZN(n436) );
  NOR2_X1 U407 ( .A1(n390), .A2(n358), .ZN(n389) );
  NOR2_X1 U408 ( .A1(n394), .A2(n392), .ZN(n390) );
  XNOR2_X1 U409 ( .A(n361), .B(n493), .ZN(n526) );
  NOR2_X1 U410 ( .A1(n611), .A2(G902), .ZN(n361) );
  XNOR2_X1 U411 ( .A(G107), .B(KEYINPUT75), .ZN(n456) );
  XOR2_X1 U412 ( .A(G104), .B(G110), .Z(n457) );
  XNOR2_X1 U413 ( .A(n414), .B(KEYINPUT39), .ZN(n542) );
  NAND2_X1 U414 ( .A1(n531), .A2(n672), .ZN(n414) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n516) );
  INV_X1 U416 ( .A(KEYINPUT73), .ZN(n359) );
  XOR2_X1 U417 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n486) );
  XNOR2_X1 U418 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n485) );
  XOR2_X1 U419 ( .A(G113), .B(G104), .Z(n484) );
  XNOR2_X1 U420 ( .A(n408), .B(G131), .ZN(n459) );
  INV_X1 U421 ( .A(G134), .ZN(n408) );
  NOR2_X1 U422 ( .A1(n734), .A2(n739), .ZN(n533) );
  AND2_X1 U423 ( .A1(G953), .A2(G902), .ZN(n428) );
  XNOR2_X1 U424 ( .A(n580), .B(n579), .ZN(n590) );
  XNOR2_X1 U425 ( .A(n578), .B(KEYINPUT87), .ZN(n579) );
  OR2_X1 U426 ( .A1(n737), .A2(KEYINPUT44), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n460), .B(n357), .ZN(n406) );
  XNOR2_X1 U428 ( .A(n459), .B(n407), .ZN(n723) );
  INV_X1 U429 ( .A(KEYINPUT94), .ZN(n407) );
  INV_X1 U430 ( .A(n654), .ZN(n373) );
  NAND2_X1 U431 ( .A1(n396), .A2(n384), .ZN(n391) );
  INV_X1 U432 ( .A(n392), .ZN(n384) );
  XNOR2_X1 U433 ( .A(n439), .B(n440), .ZN(n415) );
  OR2_X1 U434 ( .A1(n702), .A2(G902), .ZN(n416) );
  XNOR2_X1 U435 ( .A(n376), .B(n497), .ZN(n499) );
  XNOR2_X1 U436 ( .A(n496), .B(n377), .ZN(n376) );
  INV_X1 U437 ( .A(KEYINPUT103), .ZN(n377) );
  XNOR2_X1 U438 ( .A(G107), .B(G116), .ZN(n498) );
  XNOR2_X1 U439 ( .A(n481), .B(n374), .ZN(n490) );
  AND2_X2 U440 ( .A1(n383), .A2(n603), .ZN(n700) );
  XNOR2_X1 U441 ( .A(n368), .B(n468), .ZN(n469) );
  XNOR2_X1 U442 ( .A(n362), .B(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U443 ( .A1(n582), .A2(n583), .ZN(n362) );
  AND2_X1 U444 ( .A1(n512), .A2(n511), .ZN(n531) );
  XNOR2_X1 U445 ( .A(n455), .B(n454), .ZN(n466) );
  NAND2_X1 U446 ( .A1(n531), .A2(n401), .ZN(n513) );
  NOR2_X1 U447 ( .A1(n587), .A2(n402), .ZN(n401) );
  INV_X1 U448 ( .A(n507), .ZN(n402) );
  INV_X1 U449 ( .A(KEYINPUT84), .ZN(n375) );
  XNOR2_X1 U450 ( .A(KEYINPUT3), .B(G113), .ZN(n382) );
  XNOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .ZN(n421) );
  AND2_X1 U452 ( .A1(n524), .A2(n523), .ZN(n525) );
  INV_X1 U453 ( .A(KEYINPUT67), .ZN(n370) );
  XNOR2_X1 U454 ( .A(n381), .B(n379), .ZN(n472) );
  XNOR2_X1 U455 ( .A(n380), .B(G119), .ZN(n379) );
  XNOR2_X1 U456 ( .A(n382), .B(G116), .ZN(n381) );
  INV_X1 U457 ( .A(KEYINPUT70), .ZN(n380) );
  XNOR2_X1 U458 ( .A(n482), .B(KEYINPUT11), .ZN(n374) );
  XNOR2_X1 U459 ( .A(G143), .B(G131), .ZN(n482) );
  XNOR2_X1 U460 ( .A(G122), .B(G146), .ZN(n483) );
  NOR2_X1 U461 ( .A1(G237), .A2(G953), .ZN(n446) );
  XNOR2_X1 U462 ( .A(n467), .B(n369), .ZN(n368) );
  INV_X1 U463 ( .A(G125), .ZN(n369) );
  XOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n468) );
  NAND2_X1 U465 ( .A1(G237), .A2(G234), .ZN(n426) );
  NOR2_X1 U466 ( .A1(n518), .A2(n656), .ZN(n560) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(G140), .ZN(n462) );
  XNOR2_X1 U468 ( .A(n723), .B(n406), .ZN(n461) );
  NAND2_X1 U469 ( .A1(n356), .A2(n373), .ZN(n372) );
  AND2_X1 U470 ( .A1(n721), .A2(n544), .ZN(n596) );
  NOR2_X1 U471 ( .A1(n522), .A2(n521), .ZN(n538) );
  AND2_X1 U472 ( .A1(n554), .A2(n400), .ZN(n520) );
  AND2_X1 U473 ( .A1(n394), .A2(n479), .ZN(n387) );
  XNOR2_X1 U474 ( .A(n437), .B(n724), .ZN(n702) );
  XNOR2_X1 U475 ( .A(n500), .B(n378), .ZN(n605) );
  XNOR2_X1 U476 ( .A(n501), .B(n494), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n612), .B(KEYINPUT59), .ZN(n613) );
  XNOR2_X1 U478 ( .A(KEYINPUT89), .B(n608), .ZN(n705) );
  XNOR2_X1 U479 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n367) );
  INV_X1 U480 ( .A(KEYINPUT40), .ZN(n412) );
  AND2_X1 U481 ( .A1(n403), .A2(n556), .ZN(n651) );
  XNOR2_X1 U482 ( .A(n405), .B(n404), .ZN(n403) );
  XNOR2_X1 U483 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n404) );
  NAND2_X1 U484 ( .A1(n538), .A2(n507), .ZN(n405) );
  XNOR2_X1 U485 ( .A(n589), .B(KEYINPUT35), .ZN(n737) );
  NOR2_X1 U486 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U487 ( .A1(n503), .A2(n527), .ZN(n648) );
  NOR2_X1 U488 ( .A1(n503), .A2(n527), .ZN(n645) );
  INV_X1 U489 ( .A(n513), .ZN(n640) );
  AND2_X1 U490 ( .A1(G210), .A2(n480), .ZN(n353) );
  XOR2_X1 U491 ( .A(G128), .B(G146), .Z(n354) );
  XOR2_X1 U492 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n355) );
  AND2_X1 U493 ( .A1(n600), .A2(KEYINPUT2), .ZN(n356) );
  AND2_X1 U494 ( .A1(G227), .A2(n727), .ZN(n357) );
  NOR2_X1 U495 ( .A1(n671), .A2(KEYINPUT19), .ZN(n358) );
  XNOR2_X1 U496 ( .A(n421), .B(KEYINPUT90), .ZN(n604) );
  INV_X1 U497 ( .A(n604), .ZN(n398) );
  XNOR2_X2 U498 ( .A(n494), .B(n443), .ZN(n722) );
  XNOR2_X2 U499 ( .A(n442), .B(G143), .ZN(n494) );
  NOR2_X1 U500 ( .A1(n632), .A2(n644), .ZN(n564) );
  NAND2_X1 U501 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U502 ( .A1(n597), .A2(n599), .ZN(n603) );
  NAND2_X1 U503 ( .A1(n504), .A2(n642), .ZN(n360) );
  NOR2_X2 U504 ( .A1(n598), .A2(n654), .ZN(n721) );
  NAND2_X1 U505 ( .A1(n559), .A2(n553), .ZN(n363) );
  INV_X1 U506 ( .A(n557), .ZN(n365) );
  NAND2_X1 U507 ( .A1(n366), .A2(n592), .ZN(n593) );
  XNOR2_X2 U508 ( .A(n518), .B(KEYINPUT1), .ZN(n655) );
  XNOR2_X2 U509 ( .A(n464), .B(G469), .ZN(n518) );
  NAND2_X1 U510 ( .A1(n700), .A2(G475), .ZN(n614) );
  NOR2_X1 U511 ( .A1(n549), .A2(n548), .ZN(n551) );
  AND2_X1 U512 ( .A1(n565), .A2(n419), .ZN(n504) );
  NOR2_X1 U513 ( .A1(n598), .A2(n372), .ZN(n601) );
  XNOR2_X1 U514 ( .A(n537), .B(n536), .ZN(n598) );
  INV_X1 U515 ( .A(n396), .ZN(n393) );
  XNOR2_X1 U516 ( .A(n676), .B(n375), .ZN(n565) );
  NAND2_X1 U517 ( .A1(n603), .A2(n602), .ZN(n689) );
  NAND2_X1 U518 ( .A1(n393), .A2(n387), .ZN(n386) );
  NOR2_X1 U519 ( .A1(n477), .A2(n398), .ZN(n395) );
  XNOR2_X1 U520 ( .A(n470), .B(n715), .ZN(n418) );
  INV_X1 U521 ( .A(n573), .ZN(n663) );
  INV_X1 U522 ( .A(n554), .ZN(n583) );
  INV_X1 U523 ( .A(n519), .ZN(n400) );
  XNOR2_X1 U524 ( .A(n573), .B(KEYINPUT6), .ZN(n554) );
  XNOR2_X1 U525 ( .A(n435), .B(n409), .ZN(n437) );
  XNOR2_X1 U526 ( .A(n411), .B(n410), .ZN(n409) );
  XNOR2_X1 U527 ( .A(n355), .B(n433), .ZN(n410) );
  XNOR2_X1 U528 ( .A(n432), .B(n354), .ZN(n411) );
  NAND2_X1 U529 ( .A1(n542), .A2(n645), .ZN(n413) );
  XNOR2_X2 U530 ( .A(n415), .B(n416), .ZN(n659) );
  NAND2_X1 U531 ( .A1(n596), .A2(n417), .ZN(n597) );
  NAND2_X1 U532 ( .A1(n601), .A2(n417), .ZN(n602) );
  NAND2_X1 U533 ( .A1(n417), .A2(n727), .ZN(n712) );
  XNOR2_X2 U534 ( .A(n595), .B(KEYINPUT45), .ZN(n417) );
  XNOR2_X2 U535 ( .A(n458), .B(n713), .ZN(n471) );
  XNOR2_X2 U536 ( .A(n722), .B(n445), .ZN(n458) );
  XNOR2_X1 U537 ( .A(n607), .B(n606), .ZN(n609) );
  XNOR2_X1 U538 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U539 ( .A(n453), .B(G472), .ZN(n573) );
  NAND2_X1 U540 ( .A1(n700), .A2(G478), .ZN(n607) );
  XOR2_X1 U541 ( .A(KEYINPUT66), .B(KEYINPUT47), .Z(n419) );
  XNOR2_X1 U542 ( .A(n447), .B(n353), .ZN(n451) );
  INV_X1 U543 ( .A(KEYINPUT48), .ZN(n536) );
  XNOR2_X1 U544 ( .A(n469), .B(KEYINPUT79), .ZN(n470) );
  XNOR2_X1 U545 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U546 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n454) );
  XNOR2_X1 U547 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U548 ( .A(n702), .B(n701), .ZN(n703) );
  XOR2_X1 U549 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n423) );
  NAND2_X1 U550 ( .A1(n604), .A2(G234), .ZN(n422) );
  XNOR2_X1 U551 ( .A(n423), .B(n422), .ZN(n438) );
  NAND2_X1 U552 ( .A1(G221), .A2(n438), .ZN(n425) );
  XOR2_X1 U553 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n424) );
  XNOR2_X1 U554 ( .A(n425), .B(n424), .ZN(n660) );
  XOR2_X1 U555 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U556 ( .A(n427), .B(n426), .ZN(n429) );
  NAND2_X1 U557 ( .A1(G952), .A2(n429), .ZN(n684) );
  NOR2_X1 U558 ( .A1(G953), .A2(n684), .ZN(n547) );
  NAND2_X1 U559 ( .A1(n429), .A2(n428), .ZN(n545) );
  XNOR2_X1 U560 ( .A(KEYINPUT108), .B(n545), .ZN(n430) );
  NOR2_X1 U561 ( .A1(G900), .A2(n430), .ZN(n431) );
  NOR2_X1 U562 ( .A1(n547), .A2(n431), .ZN(n509) );
  XNOR2_X1 U563 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n440) );
  XOR2_X1 U564 ( .A(G119), .B(G110), .Z(n432) );
  XNOR2_X1 U565 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n433) );
  NAND2_X1 U566 ( .A1(G234), .A2(n727), .ZN(n434) );
  XOR2_X1 U567 ( .A(KEYINPUT8), .B(n434), .Z(n495) );
  NAND2_X1 U568 ( .A1(G221), .A2(n495), .ZN(n435) );
  XNOR2_X1 U569 ( .A(n460), .B(n481), .ZN(n724) );
  NAND2_X1 U570 ( .A1(G217), .A2(n438), .ZN(n439) );
  NOR2_X1 U571 ( .A1(n509), .A2(n659), .ZN(n441) );
  NAND2_X1 U572 ( .A1(n660), .A2(n441), .ZN(n519) );
  XNOR2_X2 U573 ( .A(G128), .B(KEYINPUT81), .ZN(n442) );
  INV_X1 U574 ( .A(n472), .ZN(n447) );
  XNOR2_X1 U575 ( .A(n446), .B(KEYINPUT76), .ZN(n480) );
  XOR2_X1 U576 ( .A(KEYINPUT5), .B(KEYINPUT74), .Z(n449) );
  XNOR2_X1 U577 ( .A(n459), .B(G137), .ZN(n448) );
  XNOR2_X1 U578 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U579 ( .A(n458), .B(n452), .ZN(n626) );
  NOR2_X1 U580 ( .A1(G902), .A2(n626), .ZN(n453) );
  OR2_X1 U581 ( .A1(n519), .A2(n573), .ZN(n455) );
  XNOR2_X1 U582 ( .A(n457), .B(n456), .ZN(n713) );
  XNOR2_X1 U583 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n471), .B(n463), .ZN(n693) );
  NOR2_X1 U585 ( .A1(n693), .A2(G902), .ZN(n464) );
  INV_X1 U586 ( .A(n518), .ZN(n465) );
  NAND2_X1 U587 ( .A1(n466), .A2(n465), .ZN(n529) );
  NAND2_X1 U588 ( .A1(G224), .A2(n727), .ZN(n467) );
  XNOR2_X1 U589 ( .A(G122), .B(KEYINPUT16), .ZN(n473) );
  XNOR2_X1 U590 ( .A(n473), .B(n472), .ZN(n715) );
  XOR2_X1 U591 ( .A(KEYINPUT92), .B(KEYINPUT82), .Z(n475) );
  NAND2_X1 U592 ( .A1(G210), .A2(n478), .ZN(n474) );
  XNOR2_X1 U593 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U594 ( .A(KEYINPUT91), .B(n476), .Z(n477) );
  NAND2_X1 U595 ( .A1(G214), .A2(n478), .ZN(n671) );
  INV_X1 U596 ( .A(KEYINPUT19), .ZN(n479) );
  NOR2_X2 U597 ( .A1(n529), .A2(n549), .ZN(n642) );
  NAND2_X1 U598 ( .A1(n480), .A2(G214), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n484), .B(n483), .ZN(n488) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U601 ( .A(n488), .B(n487), .Z(n489) );
  XNOR2_X1 U602 ( .A(n489), .B(n490), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n492), .B(n491), .ZN(n611) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(G475), .ZN(n493) );
  INV_X1 U605 ( .A(n526), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n495), .A2(G217), .ZN(n501) );
  XOR2_X1 U607 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n497) );
  XNOR2_X1 U608 ( .A(G122), .B(G134), .ZN(n496) );
  XNOR2_X1 U609 ( .A(n499), .B(n498), .ZN(n500) );
  NOR2_X1 U610 ( .A1(G902), .A2(n605), .ZN(n502) );
  XOR2_X1 U611 ( .A(G478), .B(n502), .Z(n527) );
  NOR2_X1 U612 ( .A1(n645), .A2(n648), .ZN(n676) );
  INV_X1 U613 ( .A(n676), .ZN(n505) );
  NAND2_X1 U614 ( .A1(n642), .A2(n505), .ZN(n506) );
  NAND2_X1 U615 ( .A1(n506), .A2(KEYINPUT47), .ZN(n514) );
  NAND2_X1 U616 ( .A1(n527), .A2(n526), .ZN(n587) );
  NAND2_X1 U617 ( .A1(n660), .A2(n659), .ZN(n656) );
  XOR2_X1 U618 ( .A(KEYINPUT110), .B(n560), .Z(n508) );
  NOR2_X1 U619 ( .A1(n509), .A2(n508), .ZN(n512) );
  NAND2_X1 U620 ( .A1(n663), .A2(n671), .ZN(n510) );
  XOR2_X1 U621 ( .A(KEYINPUT30), .B(n510), .Z(n511) );
  AND2_X1 U622 ( .A1(n514), .A2(n513), .ZN(n515) );
  AND2_X1 U623 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U624 ( .A(n517), .B(KEYINPUT72), .ZN(n524) );
  INV_X1 U625 ( .A(n645), .ZN(n522) );
  NAND2_X1 U626 ( .A1(n520), .A2(n671), .ZN(n521) );
  INV_X1 U627 ( .A(n651), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n525), .B(KEYINPUT69), .ZN(n535) );
  NAND2_X1 U629 ( .A1(n672), .A2(n671), .ZN(n675) );
  NOR2_X1 U630 ( .A1(n527), .A2(n526), .ZN(n552) );
  INV_X1 U631 ( .A(n552), .ZN(n674) );
  NOR2_X1 U632 ( .A1(n675), .A2(n674), .ZN(n528) );
  XNOR2_X1 U633 ( .A(n528), .B(KEYINPUT41), .ZN(n685) );
  NOR2_X1 U634 ( .A1(n685), .A2(n529), .ZN(n530) );
  XOR2_X1 U635 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n532) );
  XNOR2_X1 U636 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X1 U637 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n538), .A2(n655), .ZN(n539) );
  XNOR2_X1 U639 ( .A(n539), .B(KEYINPUT109), .ZN(n540) );
  XNOR2_X1 U640 ( .A(n540), .B(KEYINPUT43), .ZN(n541) );
  NOR2_X1 U641 ( .A1(n507), .A2(n541), .ZN(n654) );
  INV_X1 U642 ( .A(KEYINPUT83), .ZN(n543) );
  NAND2_X1 U643 ( .A1(n542), .A2(n648), .ZN(n720) );
  AND2_X1 U644 ( .A1(n543), .A2(n720), .ZN(n544) );
  NOR2_X1 U645 ( .A1(G898), .A2(n545), .ZN(n546) );
  NOR2_X1 U646 ( .A1(n547), .A2(n546), .ZN(n548) );
  INV_X1 U647 ( .A(KEYINPUT0), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n551), .B(n550), .ZN(n562) );
  INV_X1 U649 ( .A(n562), .ZN(n559) );
  AND2_X1 U650 ( .A1(n552), .A2(n660), .ZN(n553) );
  XNOR2_X1 U651 ( .A(n555), .B(KEYINPUT85), .ZN(n557) );
  INV_X1 U652 ( .A(n655), .ZN(n556) );
  NOR2_X1 U653 ( .A1(n655), .A2(n656), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n663), .A2(n581), .ZN(n666) );
  NOR2_X1 U655 ( .A1(n562), .A2(n666), .ZN(n563) );
  XOR2_X1 U656 ( .A(KEYINPUT31), .B(n563), .Z(n644) );
  XNOR2_X1 U657 ( .A(n564), .B(KEYINPUT99), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n420), .B(KEYINPUT104), .ZN(n567) );
  XNOR2_X1 U659 ( .A(n568), .B(KEYINPUT106), .ZN(n594) );
  INV_X1 U660 ( .A(n659), .ZN(n574) );
  NAND2_X1 U661 ( .A1(n574), .A2(n583), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n655), .A2(n569), .ZN(n570) );
  XOR2_X1 U663 ( .A(KEYINPUT80), .B(n570), .Z(n571) );
  NOR2_X1 U664 ( .A1(n576), .A2(n571), .ZN(n572) );
  XOR2_X1 U665 ( .A(KEYINPUT32), .B(n572), .Z(n738) );
  NAND2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U667 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n655), .A2(n577), .ZN(n637) );
  NAND2_X1 U669 ( .A1(n738), .A2(n637), .ZN(n580) );
  INV_X1 U670 ( .A(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n591), .A2(KEYINPUT86), .ZN(n578) );
  INV_X1 U672 ( .A(n559), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n581), .B(KEYINPUT107), .ZN(n582) );
  NOR2_X1 U674 ( .A1(n584), .A2(n686), .ZN(n586) );
  XNOR2_X1 U675 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n585) );
  XNOR2_X1 U676 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U677 ( .A1(n590), .A2(n737), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U679 ( .A(KEYINPUT2), .ZN(n599) );
  XOR2_X1 U680 ( .A(n720), .B(KEYINPUT83), .Z(n600) );
  INV_X1 U681 ( .A(n605), .ZN(n606) );
  NOR2_X1 U682 ( .A1(G952), .A2(n727), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n705), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT122), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n615), .A2(n705), .ZN(n617) );
  INV_X1 U687 ( .A(KEYINPUT60), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(G60) );
  NAND2_X1 U689 ( .A1(n700), .A2(G210), .ZN(n621) );
  XOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n618) );
  XNOR2_X1 U691 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n622), .A2(n705), .ZN(n624) );
  INV_X1 U694 ( .A(KEYINPUT56), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(G51) );
  NAND2_X1 U696 ( .A1(n700), .A2(G472), .ZN(n628) );
  XOR2_X1 U697 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n625) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n629), .A2(n705), .ZN(n631) );
  XNOR2_X1 U700 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(G57) );
  NAND2_X1 U702 ( .A1(n632), .A2(n645), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n633), .B(G104), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n635) );
  NAND2_X1 U705 ( .A1(n632), .A2(n648), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(G107), .B(n636), .ZN(G9) );
  XNOR2_X1 U708 ( .A(G110), .B(n637), .ZN(G12) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U710 ( .A1(n648), .A2(n642), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n640), .Z(n641) );
  XNOR2_X1 U713 ( .A(KEYINPUT116), .B(n641), .ZN(G45) );
  NAND2_X1 U714 ( .A1(n642), .A2(n645), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(G146), .ZN(G48) );
  XOR2_X1 U716 ( .A(G113), .B(KEYINPUT117), .Z(n647) );
  BUF_X1 U717 ( .A(n644), .Z(n649) );
  NAND2_X1 U718 ( .A1(n649), .A2(n645), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(G116), .ZN(G18) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT37), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(KEYINPUT118), .ZN(n653) );
  XNOR2_X1 U724 ( .A(G125), .B(n653), .ZN(G27) );
  XNOR2_X1 U725 ( .A(G134), .B(n720), .ZN(G36) );
  XOR2_X1 U726 ( .A(G140), .B(n654), .Z(G42) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U728 ( .A(KEYINPUT50), .B(n657), .Z(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT119), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U731 ( .A(KEYINPUT49), .B(n661), .Z(n662) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(KEYINPUT51), .B(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n685), .A2(n669), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT120), .ZN(n681) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n686), .A2(n679), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U744 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U749 ( .A1(n691), .A2(G953), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n692), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U751 ( .A(n705), .ZN(n699) );
  XNOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n693), .B(KEYINPUT57), .ZN(n694) );
  XNOR2_X1 U754 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U755 ( .A1(n700), .A2(G469), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n699), .A2(n698), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n700), .A2(G217), .ZN(n704) );
  INV_X1 U759 ( .A(KEYINPUT124), .ZN(n701) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U761 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U763 ( .A1(G224), .A2(G953), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n708), .B(KEYINPUT126), .ZN(n709) );
  XNOR2_X1 U765 ( .A(KEYINPUT61), .B(n709), .ZN(n710) );
  NAND2_X1 U766 ( .A1(n710), .A2(G898), .ZN(n711) );
  NAND2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n719) );
  XOR2_X1 U768 ( .A(G101), .B(n713), .Z(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n717) );
  NOR2_X1 U770 ( .A1(G898), .A2(n727), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(G69) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n722), .B(n723), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n725), .B(n724), .ZN(n729) );
  XNOR2_X1 U776 ( .A(n726), .B(n729), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n733) );
  XNOR2_X1 U778 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(G72) );
  XOR2_X1 U782 ( .A(n734), .B(G137), .Z(G39) );
  XNOR2_X1 U783 ( .A(n735), .B(G101), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n736), .B(KEYINPUT115), .ZN(G3) );
  XNOR2_X1 U785 ( .A(G122), .B(n737), .ZN(G24) );
  XNOR2_X1 U786 ( .A(G119), .B(n738), .ZN(G21) );
  XNOR2_X1 U787 ( .A(G131), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U788 ( .A(n740), .B(n739), .ZN(G33) );
endmodule

