//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT67), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n463), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n461), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G137), .A4(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n470), .A2(new_n479), .ZN(G160));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n473), .A2(new_n481), .A3(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n473), .B2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n473), .A2(new_n461), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n485), .A2(G124), .B1(G136), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT4), .A4(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n461), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n464), .A2(G2104), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT67), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n461), .A2(G138), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT4), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n492), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n466), .B2(new_n467), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n461), .B1(new_n497), .B2(new_n498), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n518), .ZN(G164));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n521), .B2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(KEYINPUT71), .A3(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(new_n524), .B1(KEYINPUT5), .B2(new_n521), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(G543), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n528), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  AND2_X1   g111(.A1(new_n525), .A2(new_n529), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  INV_X1    g113(.A(new_n533), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n538), .A2(new_n544), .ZN(G168));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n530), .A2(new_n546), .B1(new_n547), .B2(new_n533), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(KEYINPUT72), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(KEYINPUT72), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n527), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n527), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT74), .B(G43), .Z(new_n560));
  OAI22_X1  g135(.A1(new_n530), .A2(new_n559), .B1(new_n533), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  NAND3_X1  g143(.A1(new_n529), .A2(G53), .A3(G543), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n537), .A2(G91), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n527), .C2(new_n572), .ZN(G299));
  AND2_X1   g148(.A1(new_n554), .A2(new_n555), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  NAND3_X1  g150(.A1(new_n529), .A2(G49), .A3(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n537), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n527), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n530), .A2(new_n584), .B1(new_n585), .B2(new_n533), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n527), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n530), .A2(new_n591), .B1(new_n592), .B2(new_n533), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n537), .A2(new_n596), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n530), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n539), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n527), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  XOR2_X1   g183(.A(G284), .B(KEYINPUT76), .Z(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  INV_X1    g189(.A(new_n562), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n606), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n605), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g194(.A1(new_n485), .A2(G123), .B1(G135), .B2(new_n487), .ZN(new_n620));
  NOR2_X1   g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT77), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n507), .A2(new_n477), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT13), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT79), .B(G2443), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT80), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(G14), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT82), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n648), .ZN(new_n653));
  INV_X1    g228(.A(new_n647), .ZN(new_n654));
  OR3_X1    g229(.A1(new_n650), .A2(new_n654), .A3(new_n651), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2100), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT84), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G21), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G168), .B2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT93), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1966), .ZN(new_n688));
  NAND2_X1  g263(.A1(G299), .A2(G16), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n691));
  INV_X1    g266(.A(G20), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G1956), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT26), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n485), .B2(G129), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n477), .A2(G105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n487), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G32), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT27), .B(G1996), .Z(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G35), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G162), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT29), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n696), .B1(new_n703), .B2(new_n704), .C1(new_n708), .C2(G2090), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n487), .A2(G139), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n477), .A2(G103), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  AOI22_X1  g287(.A1(new_n507), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT90), .Z(new_n714));
  OAI211_X1 g289(.A(new_n710), .B(new_n712), .C1(new_n714), .C2(new_n461), .ZN(new_n715));
  MUX2_X1   g290(.A(G33), .B(new_n715), .S(G29), .Z(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G2072), .Z(new_n717));
  NAND2_X1  g292(.A1(G160), .A2(G29), .ZN(new_n718));
  AND2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NOR2_X1   g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n705), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(KEYINPUT91), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n705), .A2(KEYINPUT96), .A3(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n705), .ZN(new_n729));
  AOI21_X1  g304(.A(KEYINPUT96), .B1(new_n705), .B2(G27), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n717), .B(new_n727), .C1(G2078), .C2(new_n731), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n709), .B(new_n732), .C1(G29), .C2(new_n624), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT94), .B1(G5), .B2(G16), .ZN(new_n734));
  OR3_X1    g309(.A1(KEYINPUT94), .A2(G5), .A3(G16), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(G301), .C2(new_n684), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT95), .Z(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G26), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G140), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n744));
  INV_X1    g319(.A(G128), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n742), .B(new_n744), .C1(new_n484), .C2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n705), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n741), .B(new_n748), .S(KEYINPUT28), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n684), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n562), .B2(new_n684), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1341), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT31), .B(G11), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n731), .A2(G2078), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n684), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n604), .B2(new_n684), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(G28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(G28), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n762), .A2(new_n763), .A3(new_n705), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n755), .A2(new_n756), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n750), .B(new_n765), .C1(new_n703), .C2(new_n704), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n733), .A2(new_n739), .A3(new_n740), .A4(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n705), .A2(G25), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n485), .A2(G119), .B1(G131), .B2(new_n487), .ZN(new_n770));
  OR2_X1    g345(.A1(G95), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT85), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n705), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT86), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT35), .B(G1991), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n684), .A2(G24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n594), .B2(new_n684), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT87), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n684), .A2(G23), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n580), .B2(new_n684), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT88), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT33), .B(G1976), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G22), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G166), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1971), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n684), .A2(G6), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n587), .B2(new_n684), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT32), .B(G1981), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n788), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n779), .B(new_n783), .C1(new_n798), .C2(KEYINPUT34), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT89), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n688), .B(new_n768), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n708), .A2(G2090), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n724), .A2(new_n725), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n805), .A2(new_n807), .A3(new_n809), .ZN(G311));
  INV_X1    g385(.A(new_n804), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n767), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n807), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n813), .A2(new_n814), .A3(new_n808), .A4(new_n688), .ZN(G150));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n530), .A2(new_n816), .B1(new_n817), .B2(new_n533), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n525), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n527), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n604), .A2(G559), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT38), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n822), .B(KEYINPUT98), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n615), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(G860), .ZN(G145));
  NOR2_X1   g407(.A1(new_n501), .A2(new_n510), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n746), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n702), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n715), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n774), .B(new_n627), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n838));
  INV_X1    g413(.A(G106), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n461), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n487), .A2(G142), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n840), .B(new_n841), .C1(new_n485), .C2(G130), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n836), .B(new_n843), .Z(new_n844));
  XNOR2_X1  g419(.A(G160), .B(KEYINPUT99), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n624), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n836), .A2(new_n850), .A3(new_n843), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n847), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n848), .B(new_n849), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g430(.A1(new_n604), .A2(G299), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT102), .B1(new_n604), .B2(G299), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n604), .A2(G299), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n860), .B1(KEYINPUT41), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n830), .B(new_n617), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  XNOR2_X1  g444(.A(G303), .B(new_n594), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G305), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n580), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n873), .A3(KEYINPUT103), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n823), .A2(G868), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(G295));
  INV_X1    g457(.A(new_n880), .ZN(G331));
  INV_X1    g458(.A(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n867), .A2(new_n859), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n858), .B2(new_n859), .ZN(new_n886));
  XNOR2_X1  g461(.A(G168), .B(KEYINPUT105), .ZN(new_n887));
  NAND2_X1  g462(.A1(G301), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(G171), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n830), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n888), .A2(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(new_n830), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(KEYINPUT107), .A3(new_n897), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n886), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n891), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n867), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n884), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n864), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n893), .A2(new_n900), .A3(new_n894), .A4(new_n901), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n872), .B(new_n908), .C1(new_n909), .C2(new_n867), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n849), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n895), .A2(new_n902), .A3(new_n863), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n872), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n911), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n906), .A2(new_n912), .A3(new_n849), .A4(new_n910), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n915), .B2(new_n911), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(KEYINPUT44), .B2(new_n921), .ZN(G397));
  INV_X1    g497(.A(G8), .ZN(new_n923));
  INV_X1    g498(.A(G40), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n470), .A2(new_n479), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n514), .B2(new_n517), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n583), .A2(new_n586), .A3(G1981), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT49), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n932));
  INV_X1    g507(.A(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n934), .A3(new_n927), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n936), .A2(G1976), .A3(G288), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n927), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(G303), .A2(G8), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT55), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n472), .A2(new_n475), .B1(G101), .B2(new_n477), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n507), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n943));
  OAI211_X1 g518(.A(G40), .B(new_n942), .C1(new_n943), .C2(new_n461), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n511), .A2(new_n945), .A3(new_n518), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT108), .B(G1384), .ZN(new_n949));
  AOI211_X1 g524(.A(new_n947), .B(new_n949), .C1(new_n514), .C2(new_n517), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G1971), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(KEYINPUT50), .ZN(new_n953));
  INV_X1    g528(.A(G2090), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n944), .B1(new_n955), .B2(new_n926), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(G8), .B(new_n941), .C1(new_n952), .C2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n577), .A2(new_n578), .A3(G1976), .A4(new_n579), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n945), .B1(new_n501), .B2(new_n510), .ZN(new_n960));
  OAI211_X1 g535(.A(G8), .B(new_n959), .C1(new_n944), .C2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n580), .A2(G1976), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT110), .B1(new_n961), .B2(KEYINPUT52), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n961), .A2(new_n963), .A3(KEYINPUT52), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n967), .B(new_n935), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n958), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(G8), .B1(new_n952), .B2(new_n957), .ZN(new_n972));
  INV_X1    g547(.A(new_n941), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT63), .A3(new_n958), .ZN(new_n975));
  INV_X1    g550(.A(G1966), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n945), .A4(new_n518), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n925), .B1(KEYINPUT45), .B2(new_n926), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n953), .A2(new_n725), .A3(new_n956), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n508), .B1(new_n505), .B2(new_n506), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n496), .B(new_n500), .C1(new_n984), .C2(KEYINPUT4), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n985), .B2(new_n945), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n944), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n977), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT112), .A3(new_n976), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n982), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT113), .A3(G8), .A4(G168), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(G8), .A3(G168), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n970), .B(new_n975), .C1(new_n991), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n991), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n970), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n968), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n962), .A2(new_n966), .A3(new_n964), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(KEYINPUT111), .A3(new_n935), .A4(new_n967), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n948), .A2(new_n951), .ZN(new_n1004));
  INV_X1    g579(.A(G1971), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n511), .A2(new_n955), .A3(new_n945), .A4(new_n518), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n925), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n923), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n958), .B1(new_n1011), .B2(new_n941), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1003), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT63), .B1(new_n996), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n938), .B(new_n971), .C1(new_n995), .C2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G168), .A2(new_n923), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT112), .B1(new_n988), .B2(new_n976), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n981), .B(G1966), .C1(new_n987), .C2(new_n977), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n953), .A2(new_n725), .A3(new_n956), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1017), .B(new_n1020), .C1(new_n1024), .C2(new_n923), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n990), .A2(G8), .A3(G286), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1019), .C1(new_n990), .C2(G286), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(new_n1027), .A3(KEYINPUT120), .A4(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G171), .B(KEYINPUT54), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n953), .A2(new_n956), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n738), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G2078), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1035), .B1(new_n988), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1035), .B(KEYINPUT121), .C1(new_n988), .C2(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1036), .B1(new_n1004), .B2(G2078), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n958), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n944), .B(new_n950), .C1(new_n946), .C2(new_n947), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1047), .A2(G1971), .B1(G2090), .B2(new_n1009), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n941), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(KEYINPUT124), .A3(new_n998), .A4(new_n1002), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1035), .B(KEYINPUT122), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n951), .B(new_n1037), .C1(new_n1056), .C2(new_n942), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n949), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(KEYINPUT45), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1057), .A2(new_n470), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(G40), .C1(KEYINPUT123), .C2(new_n479), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1033), .A2(new_n1055), .A3(new_n1044), .A4(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1032), .A2(new_n1054), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n925), .A2(new_n926), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT116), .B(G1341), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT58), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1996), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1047), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n1071), .B2(new_n615), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n946), .A2(new_n947), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(new_n1070), .A3(new_n951), .A4(new_n925), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1068), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n562), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(KEYINPUT59), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1075), .B2(new_n562), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT117), .B(new_n615), .C1(new_n1074), .C2(new_n1068), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1009), .A2(new_n695), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(KEYINPUT115), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1073), .A2(new_n925), .A3(new_n951), .A4(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n572), .A2(new_n527), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(G91), .B2(new_n537), .ZN(new_n1090));
  NAND2_X1  g665(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1091));
  OR2_X1    g666(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1090), .A2(new_n570), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(G299), .A2(KEYINPUT114), .A3(KEYINPUT57), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1085), .A2(new_n1088), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1084), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1095), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1088), .A3(new_n1095), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1064), .B1(new_n1083), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(KEYINPUT118), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1065), .A2(G2067), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1034), .B2(new_n759), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT60), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(new_n604), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(KEYINPUT60), .B2(new_n1109), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  OR3_X1    g688(.A1(new_n1096), .A2(new_n605), .A3(new_n1109), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1101), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1015), .B1(new_n1063), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1030), .A2(new_n1118), .A3(new_n1031), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT125), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1117), .A2(new_n1125), .A3(new_n1119), .A4(new_n1122), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1116), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1059), .A2(new_n925), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1128), .A2(G1986), .A3(G290), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1128), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G1986), .A3(G290), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT109), .Z(new_n1133));
  OR2_X1    g708(.A1(new_n702), .A2(G1996), .ZN(new_n1134));
  INV_X1    g709(.A(G2067), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n746), .B(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n702), .A2(G1996), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n774), .B(new_n778), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1130), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1133), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1127), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1129), .B(KEYINPUT48), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1143), .A2(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1136), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1130), .B1(new_n702), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1130), .A2(KEYINPUT46), .A3(new_n1070), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT46), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1128), .B2(G1996), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT47), .Z(new_n1151));
  OR2_X1    g726(.A1(new_n774), .A2(new_n778), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1138), .A2(new_n1152), .B1(G2067), .B2(new_n746), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1144), .B(new_n1151), .C1(new_n1130), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1142), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1142), .A2(KEYINPUT126), .A3(new_n1154), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n1161));
  AND2_X1   g735(.A1(new_n854), .A2(new_n459), .ZN(new_n1162));
  NOR2_X1   g736(.A1(G229), .A2(G401), .ZN(new_n1163));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n661), .A3(new_n1162), .A4(new_n1163), .ZN(G225));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  NAND2_X1  g739(.A1(G225), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g740(.A(new_n1163), .ZN(new_n1167));
  AOI21_X1  g741(.A(new_n1167), .B1(new_n919), .B2(new_n920), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n1168), .A2(KEYINPUT127), .A3(new_n661), .A4(new_n1162), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1169), .ZN(G308));
endmodule


