

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U551 ( .A1(n969), .A2(n701), .ZN(n702) );
  NOR2_X1 U552 ( .A1(n627), .A2(G651), .ZN(n640) );
  NOR2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  AND2_X1 U554 ( .A1(n973), .A2(n803), .ZN(n519) );
  OR2_X1 U555 ( .A1(n757), .A2(n756), .ZN(n520) );
  XNOR2_X1 U556 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n713) );
  XNOR2_X1 U557 ( .A(n714), .B(n713), .ZN(n715) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n705) );
  XNOR2_X1 U559 ( .A(n706), .B(n705), .ZN(n711) );
  NAND2_X2 U560 ( .A1(n759), .A2(n678), .ZN(n723) );
  NAND2_X1 U561 ( .A1(G8), .A2(n723), .ZN(n752) );
  NAND2_X1 U562 ( .A1(n677), .A2(n676), .ZN(n758) );
  NOR2_X1 U563 ( .A1(n791), .A2(n519), .ZN(n792) );
  AND2_X1 U564 ( .A1(n542), .A2(n541), .ZN(n677) );
  INV_X1 U565 ( .A(G651), .ZN(n526) );
  NOR2_X1 U566 ( .A1(G543), .A2(n526), .ZN(n521) );
  XOR2_X2 U567 ( .A(KEYINPUT1), .B(n521), .Z(n639) );
  NAND2_X1 U568 ( .A1(G63), .A2(n639), .ZN(n523) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U570 ( .A1(G51), .A2(n640), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U572 ( .A(KEYINPUT6), .B(n524), .ZN(n532) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n644) );
  NAND2_X1 U574 ( .A1(n644), .A2(G89), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n525), .B(KEYINPUT4), .ZN(n528) );
  NOR2_X1 U576 ( .A1(n627), .A2(n526), .ZN(n645) );
  NAND2_X1 U577 ( .A1(G76), .A2(n645), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U579 ( .A(KEYINPUT5), .B(n529), .ZN(n530) );
  XNOR2_X1 U580 ( .A(KEYINPUT75), .B(n530), .ZN(n531) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT7), .B(n533), .Z(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U584 ( .A(G2105), .ZN(n534) );
  INV_X1 U585 ( .A(G2104), .ZN(n539) );
  NOR2_X1 U586 ( .A1(n534), .A2(n539), .ZN(n867) );
  NAND2_X1 U587 ( .A1(G113), .A2(n867), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n534), .ZN(n868) );
  NAND2_X1 U589 ( .A1(G125), .A2(n868), .ZN(n535) );
  AND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n675) );
  XOR2_X2 U591 ( .A(KEYINPUT17), .B(n537), .Z(n871) );
  NAND2_X1 U592 ( .A1(G137), .A2(n871), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n538), .B(KEYINPUT64), .ZN(n542) );
  NOR2_X2 U594 ( .A1(G2105), .A2(n539), .ZN(n872) );
  NAND2_X1 U595 ( .A1(G101), .A2(n872), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n540), .Z(n541) );
  AND2_X1 U597 ( .A1(n675), .A2(n677), .ZN(G160) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U599 ( .A1(G135), .A2(n871), .ZN(n544) );
  NAND2_X1 U600 ( .A1(G111), .A2(n867), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n868), .A2(G123), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(n545), .Z(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n872), .A2(G99), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n937) );
  XNOR2_X1 U607 ( .A(G2096), .B(n937), .ZN(n550) );
  OR2_X1 U608 ( .A1(G2100), .A2(n550), .ZN(G156) );
  XNOR2_X1 U609 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n644), .A2(G81), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT12), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G68), .A2(n645), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U614 ( .A(n555), .B(n554), .Z(n560) );
  XOR2_X1 U615 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n557) );
  NAND2_X1 U616 ( .A1(G56), .A2(n639), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U618 ( .A(KEYINPUT69), .B(n558), .ZN(n559) );
  AND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT72), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G43), .A2(n640), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n687) );
  INV_X1 U623 ( .A(G860), .ZN(n815) );
  OR2_X1 U624 ( .A1(n687), .A2(n815), .ZN(G153) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G82), .ZN(G220) );
  NAND2_X1 U627 ( .A1(G64), .A2(n639), .ZN(n565) );
  NAND2_X1 U628 ( .A1(G52), .A2(n640), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G90), .A2(n644), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G77), .A2(n645), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U634 ( .A1(n570), .A2(n569), .ZN(G171) );
  NAND2_X1 U635 ( .A1(G138), .A2(n871), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G102), .A2(n872), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G114), .A2(n867), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G126), .A2(n868), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(G164) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n808) );
  NAND2_X1 U645 ( .A1(n808), .A2(G567), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G54), .A2(n640), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G92), .A2(n644), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G79), .A2(n645), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G66), .A2(n639), .ZN(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT73), .B(n581), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT15), .ZN(n587) );
  XNOR2_X2 U657 ( .A(KEYINPUT74), .B(n587), .ZN(n959) );
  INV_X1 U658 ( .A(n959), .ZN(n885) );
  NOR2_X1 U659 ( .A1(n885), .A2(G868), .ZN(n589) );
  INV_X1 U660 ( .A(G868), .ZN(n659) );
  NOR2_X1 U661 ( .A1(n659), .A2(G301), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G91), .A2(n644), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT66), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G65), .A2(n639), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G53), .A2(n640), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G78), .A2(n645), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT67), .B(n593), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n659), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U675 ( .A1(G559), .A2(n815), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n600), .B(KEYINPUT76), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n601), .A2(n959), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT16), .B(n602), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n687), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n959), .A2(G868), .ZN(n603) );
  NOR2_X1 U681 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G86), .A2(n644), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G61), .A2(n639), .ZN(n606) );
  XNOR2_X1 U685 ( .A(n606), .B(KEYINPUT80), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G73), .A2(n645), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G48), .A2(n640), .ZN(n610) );
  XNOR2_X1 U690 ( .A(KEYINPUT81), .B(n610), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U694 ( .A1(G88), .A2(n644), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G75), .A2(n645), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U697 ( .A(KEYINPUT84), .B(n618), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G62), .A2(n639), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT83), .B(n619), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n640), .A2(G50), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(G303) );
  INV_X1 U703 ( .A(G303), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G49), .A2(n640), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n639), .A2(n626), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G60), .A2(n639), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G47), .A2(n640), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G85), .A2(n644), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G72), .A2(n645), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n636), .B(KEYINPUT65), .ZN(G290) );
  XNOR2_X1 U718 ( .A(n687), .B(KEYINPUT77), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n959), .A2(G559), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n638), .B(n637), .ZN(n814) );
  NAND2_X1 U721 ( .A1(G67), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G55), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U724 ( .A(KEYINPUT78), .B(n643), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G93), .A2(n644), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G80), .A2(n645), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U729 ( .A(KEYINPUT79), .B(n650), .ZN(n816) );
  XOR2_X1 U730 ( .A(G305), .B(n816), .Z(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n652) );
  XNOR2_X1 U732 ( .A(G288), .B(KEYINPUT86), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(G166), .B(n653), .ZN(n655) );
  INV_X1 U735 ( .A(G299), .ZN(n969) );
  XNOR2_X1 U736 ( .A(G290), .B(n969), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n657), .B(n656), .ZN(n884) );
  XNOR2_X1 U739 ( .A(n814), .B(n884), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n658), .A2(G868), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n659), .A2(n816), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G108), .A2(G120), .ZN(n666) );
  NOR2_X1 U751 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U752 ( .A1(G69), .A2(n667), .ZN(n812) );
  NAND2_X1 U753 ( .A1(n812), .A2(G567), .ZN(n672) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U756 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(G96), .A2(n670), .ZN(n813) );
  NAND2_X1 U758 ( .A1(n813), .A2(G2106), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n672), .A2(n671), .ZN(n818) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n673) );
  NOR2_X1 U761 ( .A1(n818), .A2(n673), .ZN(n811) );
  NAND2_X1 U762 ( .A1(n811), .A2(G36), .ZN(n674) );
  XOR2_X1 U763 ( .A(KEYINPUT87), .B(n674), .Z(G176) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n759) );
  AND2_X1 U765 ( .A1(n675), .A2(G40), .ZN(n676) );
  INV_X1 U766 ( .A(n758), .ZN(n678) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n679) );
  XOR2_X1 U768 ( .A(n679), .B(KEYINPUT24), .Z(n680) );
  NOR2_X1 U769 ( .A1(n752), .A2(n680), .ZN(n757) );
  INV_X1 U770 ( .A(n723), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n707), .A2(G1348), .ZN(n682) );
  NOR2_X1 U772 ( .A1(G2067), .A2(n723), .ZN(n681) );
  NOR2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n707), .A2(G1996), .ZN(n683) );
  XNOR2_X1 U775 ( .A(n683), .B(KEYINPUT26), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n723), .A2(G1341), .ZN(n684) );
  NAND2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n691), .A2(n959), .ZN(n688) );
  NAND2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U780 ( .A(KEYINPUT95), .B(n690), .Z(n693) );
  OR2_X1 U781 ( .A1(n959), .A2(n691), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n700) );
  NAND2_X1 U783 ( .A1(n707), .A2(G2072), .ZN(n695) );
  INV_X1 U784 ( .A(KEYINPUT27), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n723), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U788 ( .A(KEYINPUT94), .B(n698), .Z(n701) );
  NAND2_X1 U789 ( .A1(n969), .A2(n701), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n704) );
  XOR2_X1 U791 ( .A(n702), .B(KEYINPUT28), .Z(n703) );
  NAND2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U793 ( .A(KEYINPUT25), .B(G2078), .Z(n909) );
  NOR2_X1 U794 ( .A1(n909), .A2(n723), .ZN(n709) );
  NOR2_X1 U795 ( .A1(n707), .A2(G1961), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n717) );
  OR2_X1 U797 ( .A1(n717), .A2(G301), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n722) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n752), .ZN(n732) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n723), .ZN(n731) );
  NOR2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n712) );
  NAND2_X1 U802 ( .A1(G8), .A2(n712), .ZN(n714) );
  NOR2_X1 U803 ( .A1(G168), .A2(n715), .ZN(n716) );
  XNOR2_X1 U804 ( .A(n716), .B(KEYINPUT97), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n717), .A2(G301), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT31), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n733), .A2(G286), .ZN(n728) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n752), .ZN(n725) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U814 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U816 ( .A(n730), .B(KEYINPUT32), .ZN(n738) );
  NAND2_X1 U817 ( .A1(G8), .A2(n731), .ZN(n736) );
  INV_X1 U818 ( .A(n733), .ZN(n734) );
  NOR2_X1 U819 ( .A1(n732), .A2(n734), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n738), .A2(n737), .ZN(n751) );
  NOR2_X1 U822 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U823 ( .A1(G1971), .A2(G303), .ZN(n739) );
  NOR2_X1 U824 ( .A1(n744), .A2(n739), .ZN(n965) );
  NAND2_X1 U825 ( .A1(n751), .A2(n965), .ZN(n740) );
  NAND2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n964) );
  NAND2_X1 U827 ( .A1(n740), .A2(n964), .ZN(n741) );
  XNOR2_X1 U828 ( .A(KEYINPUT98), .B(n741), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n742), .A2(n752), .ZN(n743) );
  NOR2_X1 U830 ( .A1(KEYINPUT33), .A2(n743), .ZN(n747) );
  NAND2_X1 U831 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n745), .A2(n752), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U834 ( .A(G1981), .B(G305), .Z(n956) );
  NAND2_X1 U835 ( .A1(n748), .A2(n956), .ZN(n755) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n749) );
  NAND2_X1 U837 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n759), .A2(n758), .ZN(n803) );
  XNOR2_X1 U842 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  XNOR2_X1 U843 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n763) );
  NAND2_X1 U844 ( .A1(G116), .A2(n867), .ZN(n761) );
  NAND2_X1 U845 ( .A1(G128), .A2(n868), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U847 ( .A(n763), .B(n762), .ZN(n769) );
  NAND2_X1 U848 ( .A1(n872), .A2(G104), .ZN(n764) );
  XNOR2_X1 U849 ( .A(n764), .B(KEYINPUT88), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G140), .A2(n871), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(n767), .ZN(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U854 ( .A(KEYINPUT36), .B(n770), .ZN(n846) );
  NOR2_X1 U855 ( .A1(n801), .A2(n846), .ZN(n949) );
  NAND2_X1 U856 ( .A1(n803), .A2(n949), .ZN(n799) );
  NAND2_X1 U857 ( .A1(G105), .A2(n872), .ZN(n771) );
  XOR2_X1 U858 ( .A(KEYINPUT38), .B(n771), .Z(n776) );
  NAND2_X1 U859 ( .A1(G117), .A2(n867), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G129), .A2(n868), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U862 ( .A(KEYINPUT91), .B(n774), .Z(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n871), .A2(G141), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n878) );
  NAND2_X1 U866 ( .A1(G1996), .A2(n878), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(KEYINPUT92), .ZN(n788) );
  NAND2_X1 U868 ( .A1(G131), .A2(n871), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G119), .A2(n868), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n867), .A2(G107), .ZN(n782) );
  XOR2_X1 U872 ( .A(KEYINPUT90), .B(n782), .Z(n783) );
  NOR2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n872), .A2(G95), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n858) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n858), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n936) );
  NAND2_X1 U878 ( .A1(n936), .A2(n803), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT93), .ZN(n796) );
  INV_X1 U880 ( .A(n796), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n799), .A2(n790), .ZN(n791) );
  XNOR2_X1 U882 ( .A(G1986), .B(G290), .ZN(n973) );
  NAND2_X1 U883 ( .A1(n520), .A2(n792), .ZN(n806) );
  NOR2_X1 U884 ( .A1(G1996), .A2(n878), .ZN(n933) );
  NOR2_X1 U885 ( .A1(G1986), .A2(G290), .ZN(n793) );
  XOR2_X1 U886 ( .A(n793), .B(KEYINPUT99), .Z(n794) );
  NOR2_X1 U887 ( .A1(G1991), .A2(n858), .ZN(n940) );
  NOR2_X1 U888 ( .A1(n794), .A2(n940), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U890 ( .A1(n933), .A2(n797), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT39), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n801), .A2(n846), .ZN(n946) );
  NAND2_X1 U894 ( .A1(n802), .A2(n946), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U897 ( .A(n807), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U898 ( .A1(G2106), .A2(n808), .ZN(G217) );
  AND2_X1 U899 ( .A1(G15), .A2(G2), .ZN(n809) );
  NAND2_X1 U900 ( .A1(G661), .A2(n809), .ZN(G259) );
  NAND2_X1 U901 ( .A1(G3), .A2(G1), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(G188) );
  INV_X1 U904 ( .A(G120), .ZN(G236) );
  INV_X1 U905 ( .A(G108), .ZN(G238) );
  INV_X1 U906 ( .A(G96), .ZN(G221) );
  INV_X1 U907 ( .A(G69), .ZN(G235) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(G325) );
  INV_X1 U909 ( .A(G325), .ZN(G261) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(n816), .ZN(G145) );
  INV_X1 U912 ( .A(n818), .ZN(G319) );
  XOR2_X1 U913 ( .A(G2678), .B(KEYINPUT43), .Z(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT42), .B(G2090), .Z(n822) );
  XNOR2_X1 U917 ( .A(G2067), .B(G2072), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U919 ( .A(n824), .B(n823), .Z(n826) );
  XNOR2_X1 U920 ( .A(G2096), .B(G2100), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n826), .B(n825), .ZN(n828) );
  XOR2_X1 U922 ( .A(G2078), .B(G2084), .Z(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(G227) );
  XOR2_X1 U924 ( .A(G1976), .B(G1971), .Z(n830) );
  XNOR2_X1 U925 ( .A(G1986), .B(G1961), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U927 ( .A(n831), .B(G2474), .Z(n833) );
  XNOR2_X1 U928 ( .A(G1966), .B(G1981), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT41), .B(G1956), .Z(n835) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(G229) );
  NAND2_X1 U934 ( .A1(G124), .A2(n868), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT44), .ZN(n841) );
  NAND2_X1 U936 ( .A1(G100), .A2(n872), .ZN(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT103), .B(n839), .Z(n840) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G136), .A2(n871), .ZN(n843) );
  NAND2_X1 U940 ( .A1(G112), .A2(n867), .ZN(n842) );
  NAND2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(G162) );
  XNOR2_X1 U943 ( .A(G160), .B(n846), .ZN(n857) );
  NAND2_X1 U944 ( .A1(G139), .A2(n871), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT106), .ZN(n856) );
  NAND2_X1 U946 ( .A1(n872), .A2(G103), .ZN(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT105), .B(n848), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G115), .A2(n867), .ZN(n850) );
  NAND2_X1 U949 ( .A1(G127), .A2(n868), .ZN(n849) );
  NAND2_X1 U950 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT107), .B(n851), .ZN(n852) );
  XNOR2_X1 U952 ( .A(KEYINPUT47), .B(n852), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n927) );
  XNOR2_X1 U955 ( .A(n857), .B(n927), .ZN(n861) );
  XNOR2_X1 U956 ( .A(G164), .B(n858), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(n937), .ZN(n860) );
  XOR2_X1 U958 ( .A(n861), .B(n860), .Z(n866) );
  XOR2_X1 U959 ( .A(KEYINPUT104), .B(KEYINPUT46), .Z(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT48), .B(KEYINPUT108), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT109), .B(n864), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n882) );
  NAND2_X1 U964 ( .A1(G118), .A2(n867), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G130), .A2(n868), .ZN(n869) );
  NAND2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U967 ( .A1(G142), .A2(n871), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G106), .A2(n872), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U970 ( .A(n875), .B(KEYINPUT45), .Z(n876) );
  NOR2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n879) );
  XNOR2_X1 U972 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U973 ( .A(G162), .B(n880), .Z(n881) );
  XNOR2_X1 U974 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U975 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U976 ( .A(G286), .B(n884), .ZN(n889) );
  XOR2_X1 U977 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n887) );
  XNOR2_X1 U978 ( .A(G171), .B(n885), .ZN(n886) );
  XNOR2_X1 U979 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U981 ( .A(n890), .B(n687), .Z(n891) );
  NOR2_X1 U982 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U983 ( .A(KEYINPUT100), .B(G2446), .Z(n893) );
  XNOR2_X1 U984 ( .A(G2443), .B(G2454), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U986 ( .A(n894), .B(G2451), .Z(n896) );
  XNOR2_X1 U987 ( .A(G1341), .B(G1348), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n896), .B(n895), .ZN(n900) );
  XOR2_X1 U989 ( .A(G2435), .B(G2427), .Z(n898) );
  XNOR2_X1 U990 ( .A(G2430), .B(G2438), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U992 ( .A(n900), .B(n899), .Z(n901) );
  NAND2_X1 U993 ( .A1(G14), .A2(n901), .ZN(n907) );
  NAND2_X1 U994 ( .A1(G319), .A2(n907), .ZN(n904) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n902) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U997 ( .A1(n904), .A2(n903), .ZN(n906) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(n907), .ZN(G401) );
  XNOR2_X1 U1002 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1017) );
  XOR2_X1 U1003 ( .A(G1991), .B(G25), .Z(n908) );
  NAND2_X1 U1004 ( .A1(n908), .A2(G28), .ZN(n914) );
  XNOR2_X1 U1005 ( .A(G1996), .B(G32), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n909), .B(G27), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT116), .B(n912), .Z(n913) );
  NOR2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(G33), .B(G2072), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(KEYINPUT53), .ZN(n922) );
  XOR2_X1 U1015 ( .A(G2084), .B(G34), .Z(n920) );
  XNOR2_X1 U1016 ( .A(KEYINPUT54), .B(n920), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(G35), .B(G2090), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1020 ( .A(KEYINPUT55), .B(n925), .Z(n926) );
  NOR2_X1 U1021 ( .A1(G29), .A2(n926), .ZN(n1015) );
  INV_X1 U1022 ( .A(KEYINPUT55), .ZN(n953) );
  XNOR2_X1 U1023 ( .A(KEYINPUT52), .B(KEYINPUT114), .ZN(n951) );
  XNOR2_X1 U1024 ( .A(G164), .B(G2078), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(G2072), .B(KEYINPUT113), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT50), .ZN(n945) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n934), .B(KEYINPUT51), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(KEYINPUT112), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(n951), .B(n950), .ZN(n952) );
  NAND2_X1 U1042 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1043 ( .A1(n954), .A2(G29), .ZN(n955) );
  XNOR2_X1 U1044 ( .A(n955), .B(KEYINPUT115), .ZN(n1012) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n981) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G168), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(KEYINPUT57), .B(n958), .ZN(n979) );
  XNOR2_X1 U1049 ( .A(G171), .B(G1961), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(n959), .B(G1348), .ZN(n960) );
  NAND2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G1341), .B(n687), .ZN(n962) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n976) );
  NAND2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n967) );
  AND2_X1 U1055 ( .A1(G303), .A2(G1971), .ZN(n966) );
  NOR2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1057 ( .A(KEYINPUT117), .B(n968), .Z(n971) );
  XNOR2_X1 U1058 ( .A(n969), .B(G1956), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1060 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1061 ( .A(n974), .B(KEYINPUT118), .ZN(n975) );
  NAND2_X1 U1062 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(KEYINPUT119), .B(n977), .ZN(n978) );
  NAND2_X1 U1064 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1065 ( .A1(n981), .A2(n980), .ZN(n1010) );
  XOR2_X1 U1066 ( .A(G16), .B(KEYINPUT120), .Z(n1008) );
  XOR2_X1 U1067 ( .A(G1986), .B(G24), .Z(n984) );
  XOR2_X1 U1068 ( .A(G22), .B(KEYINPUT124), .Z(n982) );
  XNOR2_X1 U1069 ( .A(n982), .B(G1971), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1071 ( .A(KEYINPUT125), .B(G1976), .Z(n985) );
  XNOR2_X1 U1072 ( .A(G23), .B(n985), .ZN(n986) );
  NOR2_X1 U1073 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1074 ( .A(KEYINPUT58), .B(n988), .Z(n1005) );
  XOR2_X1 U1075 ( .A(G1961), .B(G5), .Z(n1000) );
  XNOR2_X1 U1076 ( .A(KEYINPUT59), .B(G1348), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n989), .B(G4), .ZN(n996) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G20), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G1981), .B(G6), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT121), .B(n992), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT122), .B(n997), .Z(n998) );
  XNOR2_X1 U1086 ( .A(n998), .B(KEYINPUT60), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G21), .B(G1966), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(KEYINPUT123), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(KEYINPUT61), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1095 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1096 ( .A1(n1013), .A2(G11), .ZN(n1014) );
  NOR2_X1 U1097 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1017), .B(n1016), .ZN(G311) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

