//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT28), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT72), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n206));
  NAND4_X1  g005(.A1(new_n202), .A2(new_n206), .A3(KEYINPUT28), .A4(new_n203), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT27), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n203), .B(new_n212), .C1(new_n202), .C2(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n203), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n209), .B(new_n214), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n208), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n214), .B1(new_n219), .B2(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT71), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n221), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT73), .A3(new_n208), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n211), .A2(new_n203), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT69), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT26), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n229), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT64), .Z(new_n245));
  OR3_X1    g044(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n211), .B2(new_n203), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G169gat), .B2(G176gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n252), .A2(new_n237), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(new_n246), .A2(new_n249), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n244), .B(KEYINPUT64), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n248), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n256), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n251), .A2(new_n257), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n244), .B1(G183gat), .B2(G190gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n231), .B2(new_n247), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(KEYINPUT25), .A3(new_n254), .A4(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n253), .B1(new_n233), .B2(new_n235), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n267), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n243), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT77), .A2(G113gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT77), .A2(G113gat), .ZN(new_n277));
  OAI21_X1  g076(.A(G120gat), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(KEYINPUT78), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT1), .B1(new_n283), .B2(G127gat), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G134gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n284), .B(new_n286), .C1(new_n278), .C2(KEYINPUT78), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT79), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(KEYINPUT77), .A2(G113gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT77), .A2(G113gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n279), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(new_n285), .B2(G134gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n284), .A4(new_n281), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT76), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT75), .B(G134gat), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n297), .B(new_n286), .C1(new_n298), .C2(new_n285), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n283), .A2(KEYINPUT75), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n283), .A2(KEYINPUT75), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT76), .B(G127gat), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  INV_X1    g102(.A(new_n280), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n279), .A2(G113gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT80), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n288), .B2(new_n295), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n275), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G227gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n243), .A2(new_n309), .A3(new_n274), .A4(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G15gat), .B(G43gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT34), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n315), .A2(new_n319), .ZN(new_n329));
  INV_X1    g128(.A(new_n318), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI211_X1 g130(.A(KEYINPUT34), .B(new_n318), .C1(new_n315), .C2(new_n319), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n327), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n334));
  INV_X1    g133(.A(new_n319), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n243), .A2(new_n274), .B1(new_n309), .B2(new_n313), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT34), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(new_n328), .A3(new_n330), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n326), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  INV_X1    g141(.A(new_n326), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n338), .A2(new_n339), .A3(new_n334), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n341), .A2(KEYINPUT36), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT36), .B1(new_n341), .B2(new_n345), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT82), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n272), .B1(new_n263), .B2(new_n264), .ZN(new_n351));
  AOI221_X4 g150(.A(new_n224), .B1(new_n205), .B2(new_n207), .C1(new_n227), .C2(new_n221), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT73), .B1(new_n228), .B2(new_n208), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n354), .B2(new_n242), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n348), .B(new_n350), .C1(new_n355), .C2(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT29), .B1(new_n243), .B2(new_n274), .ZN(new_n357));
  INV_X1    g156(.A(new_n350), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT83), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT22), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n362), .B2(new_n363), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n365), .A2(KEYINPUT81), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n367), .A2(KEYINPUT81), .A3(new_n360), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n349), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n275), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n359), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n370), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n371), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n355), .A2(new_n350), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(G64gat), .ZN(new_n380));
  INV_X1    g179(.A(G92gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n373), .A2(new_n377), .A3(new_n382), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n378), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  XOR2_X1   g187(.A(G155gat), .B(G162gat), .Z(new_n389));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(G155gat), .B2(G162gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G141gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G148gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT85), .B(G148gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n393), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT84), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT84), .B1(new_n394), .B2(new_n400), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n391), .ZN(new_n403));
  INV_X1    g202(.A(new_n389), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n397), .B(new_n398), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n308), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n311), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n296), .A2(new_n312), .A3(new_n307), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n312), .B1(new_n296), .B2(new_n307), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n408), .B(new_n414), .C1(new_n417), .C2(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n308), .A2(new_n406), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT86), .A3(new_n412), .ZN(new_n420));
  OR3_X1    g219(.A1(new_n311), .A2(KEYINPUT86), .A3(new_n411), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n410), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(KEYINPUT5), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n405), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n412), .A2(new_n413), .B1(new_n424), .B2(new_n311), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n413), .B2(new_n417), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n409), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT0), .B(G57gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n434), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n423), .A2(new_n428), .A3(new_n433), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n386), .A2(new_n388), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT29), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n368), .B2(new_n369), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n411), .B1(new_n443), .B2(new_n398), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n405), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n370), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(new_n445), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n451), .B1(new_n444), .B2(KEYINPUT88), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(new_n448), .C1(KEYINPUT88), .C2(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n441), .B1(new_n455), .B2(G22gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n452), .A2(new_n461), .A3(new_n454), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n452), .B2(new_n454), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n456), .A2(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n466), .A2(new_n441), .A3(new_n462), .A4(new_n459), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n346), .A2(new_n347), .B1(new_n440), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n435), .A3(new_n384), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n383), .B1(new_n378), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n471), .B2(new_n378), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(KEYINPUT38), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n356), .A2(new_n359), .A3(new_n374), .A4(new_n372), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT92), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n475), .B(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n480), .A3(KEYINPUT37), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n474), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n465), .A2(new_n467), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT4), .B1(new_n314), .B2(new_n411), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n410), .B1(new_n490), .B2(new_n425), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n420), .A2(new_n421), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n409), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n491), .A2(KEYINPUT39), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n426), .A2(KEYINPUT39), .A3(new_n409), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n434), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT90), .B(new_n433), .C1(new_n491), .C2(KEYINPUT39), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT40), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n436), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n501), .B(new_n494), .C1(new_n497), .C2(new_n498), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n386), .A2(new_n388), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n489), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n469), .B1(new_n488), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n468), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n439), .A2(new_n435), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n440), .A2(new_n514), .A3(KEYINPUT35), .A4(new_n468), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G22gat), .Z(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT16), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n526), .B(KEYINPUT95), .Z(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n527), .B2(new_n523), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT96), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n528), .B(new_n531), .Z(new_n532));
  AOI21_X1  g331(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT99), .ZN(new_n534));
  XOR2_X1   g333(.A(G57gat), .B(G64gat), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(KEYINPUT99), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(new_n211), .ZN(new_n542));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(new_n362), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n544), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n547), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G43gat), .B(G50gat), .Z(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OR3_X1    g354(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n556), .A2(new_n557), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n553), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(KEYINPUT15), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n562), .A3(new_n558), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT17), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT97), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n570), .B2(new_n381), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G99gat), .B(G106gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT101), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n563), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT94), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT102), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n581), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n576), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n586), .A2(new_n587), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n565), .A2(new_n590), .A3(new_n576), .A4(new_n582), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n584), .A2(new_n595), .A3(new_n589), .A4(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n594), .A2(new_n600), .A3(new_n596), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT11), .B(G169gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G197gat), .ZN(new_n606));
  XOR2_X1   g405(.A(G113gat), .B(G141gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n565), .A2(new_n532), .A3(new_n582), .ZN(new_n610));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n585), .A2(new_n532), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT18), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n585), .B(new_n532), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n611), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT18), .A4(new_n611), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n615), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n617), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G230gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n317), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n576), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n539), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n573), .A2(new_n575), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n573), .A2(new_n575), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT103), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n576), .A2(new_n628), .A3(new_n539), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT10), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n576), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n627), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(new_n626), .A3(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G176gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT104), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT105), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648));
  AOI211_X1 g447(.A(new_n648), .B(new_n645), .C1(new_n639), .C2(new_n640), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n641), .A2(new_n644), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n624), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n552), .A2(new_n604), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n522), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n516), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g456(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n658));
  OR2_X1    g457(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n654), .A2(new_n507), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT107), .B1(new_n660), .B2(KEYINPUT106), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n662));
  INV_X1    g461(.A(new_n654), .ZN(new_n663));
  OAI21_X1  g462(.A(G8gat), .B1(new_n663), .B2(new_n506), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n660), .B2(KEYINPUT107), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n662), .B(new_n664), .C1(new_n666), .C2(new_n661), .ZN(G1325gat));
  AOI21_X1  g466(.A(G15gat), .B1(new_n654), .B2(new_n514), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n654), .A2(G15gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n346), .A2(new_n347), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n489), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  OAI21_X1  g473(.A(new_n604), .B1(new_n509), .B2(new_n520), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n604), .C1(new_n509), .C2(new_n520), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n551), .A2(new_n652), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT109), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n677), .A2(new_n682), .A3(new_n678), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n655), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n685), .A2(KEYINPUT110), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(KEYINPUT110), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(G29gat), .A3(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n675), .A2(new_n551), .A3(new_n652), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(new_n655), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n688), .A2(new_n694), .A3(new_n695), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G36gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n689), .A2(new_n700), .A3(new_n507), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n506), .B1(new_n681), .B2(new_n683), .ZN(new_n704));
  OAI221_X1 g503(.A(new_n703), .B1(new_n699), .B2(new_n701), .C1(new_n704), .C2(new_n700), .ZN(G1329gat));
  INV_X1    g504(.A(new_n670), .ZN(new_n706));
  OAI21_X1  g505(.A(G43gat), .B1(new_n680), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n689), .A2(new_n708), .A3(new_n514), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n684), .B2(new_n670), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT112), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n711), .B(new_n717), .C1(new_n712), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n680), .B2(new_n468), .ZN(new_n720));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n689), .A2(new_n721), .A3(new_n489), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(KEYINPUT48), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n468), .B1(new_n681), .B2(new_n683), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n604), .ZN(new_n731));
  INV_X1    g530(.A(new_n624), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n551), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n510), .B2(new_n521), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n516), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g537(.A1(new_n736), .A2(new_n506), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND4_X1  g542(.A1(new_n734), .A2(G71gat), .A3(new_n670), .A4(new_n735), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n736), .A2(new_n512), .A3(new_n513), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(G71gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n736), .A2(new_n468), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT114), .B(G78gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n551), .A2(new_n624), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n677), .A2(new_n735), .A3(new_n678), .A4(new_n751), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n570), .A3(new_n516), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(new_n751), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n675), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n675), .B2(new_n755), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(KEYINPUT115), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n735), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n655), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n753), .B1(new_n764), .B2(new_n570), .ZN(G1336gat));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g565(.A(G92gat), .B1(new_n752), .B2(new_n506), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n507), .A2(new_n381), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n762), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n651), .B1(new_n757), .B2(new_n758), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n381), .A3(new_n507), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n771), .A2(new_n767), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(new_n766), .ZN(G1337gat));
  INV_X1    g572(.A(G99gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n763), .A2(new_n774), .A3(new_n514), .ZN(new_n775));
  OAI21_X1  g574(.A(G99gat), .B1(new_n752), .B2(new_n706), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1338gat));
  NOR2_X1   g576(.A1(new_n468), .A2(G106gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n759), .A2(new_n735), .A3(new_n761), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  OAI21_X1  g579(.A(G106gat), .B1(new_n752), .B2(new_n468), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n770), .A2(new_n778), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(new_n781), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT116), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n783), .A2(new_n781), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n780), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1339gat));
  NOR2_X1   g589(.A1(new_n733), .A2(new_n735), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n627), .C1(new_n636), .C2(new_n638), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n644), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n634), .A2(new_n635), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n638), .B1(new_n796), .B2(new_n637), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n626), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n639), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n799), .A3(KEYINPUT55), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n795), .A2(new_n799), .A3(KEYINPUT117), .A4(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n795), .B2(new_n799), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n650), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n624), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n615), .A2(new_n621), .A3(new_n609), .A4(new_n622), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n618), .A2(new_n620), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n608), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n735), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n604), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n602), .B2(new_n603), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n804), .A2(new_n816), .A3(new_n806), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n552), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n792), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n515), .A2(new_n507), .A3(new_n516), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n732), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n821), .B(KEYINPUT118), .Z(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n277), .B2(new_n276), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(new_n732), .ZN(G1340gat));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n279), .A3(new_n735), .ZN(new_n826));
  OAI21_X1  g625(.A(G120gat), .B1(new_n821), .B2(new_n651), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  NOR2_X1   g627(.A1(new_n821), .A2(new_n552), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(new_n285), .ZN(G1342gat));
  NOR3_X1   g629(.A1(new_n821), .A2(new_n298), .A3(new_n731), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n821), .B2(new_n731), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n489), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n670), .A2(new_n516), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n507), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n651), .B2(new_n812), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n735), .A2(new_n845), .A3(new_n813), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n807), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n731), .ZN(new_n848));
  INV_X1    g647(.A(new_n817), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n552), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n792), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n843), .B1(new_n852), .B2(new_n489), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n842), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n393), .B1(new_n854), .B2(new_n624), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n468), .B1(new_n792), .B2(new_n818), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n732), .A2(G141gat), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n506), .A3(new_n839), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT120), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n839), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n507), .B1(new_n862), .B2(KEYINPUT121), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(KEYINPUT121), .B2(new_n862), .ZN(new_n864));
  INV_X1    g663(.A(new_n857), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n860), .B1(new_n855), .B2(new_n866), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n854), .A2(new_n735), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n395), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT122), .B1(new_n848), .B2(new_n849), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(new_n817), .C1(new_n847), .C2(new_n731), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(new_n874), .A3(new_n551), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n843), .B(new_n489), .C1(new_n875), .C2(new_n791), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n735), .A3(new_n877), .A4(new_n841), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G148gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n871), .B1(new_n879), .B2(KEYINPUT59), .ZN(new_n880));
  AOI211_X1 g679(.A(KEYINPUT123), .B(new_n869), .C1(new_n878), .C2(G148gat), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n864), .A2(new_n395), .A3(new_n651), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n864), .A2(new_n552), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n854), .A2(new_n551), .ZN(new_n886));
  MUX2_X1   g685(.A(new_n885), .B(new_n886), .S(G155gat), .Z(G1346gat));
  NOR2_X1   g686(.A1(new_n864), .A2(new_n731), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n854), .A2(new_n604), .ZN(new_n889));
  MUX2_X1   g688(.A(new_n888), .B(new_n889), .S(G162gat), .Z(G1347gat));
  NOR2_X1   g689(.A1(new_n655), .A2(new_n506), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n515), .B(new_n892), .C1(new_n792), .C2(new_n818), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n624), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n735), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(G176gat), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT124), .B(G176gat), .Z(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n896), .B2(new_n899), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n551), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n211), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n202), .B2(new_n901), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g703(.A1(new_n893), .A2(new_n604), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(new_n203), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT61), .B(G190gat), .Z(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n905), .B2(new_n908), .ZN(G1351gat));
  NAND2_X1  g708(.A1(new_n850), .A2(new_n873), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n848), .A2(KEYINPUT122), .A3(new_n849), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n552), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n792), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n913), .A2(new_n489), .B1(KEYINPUT57), .B2(new_n837), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n892), .A2(new_n670), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n732), .ZN(new_n917));
  INV_X1    g716(.A(new_n915), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n837), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n624), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n917), .A2(new_n921), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n735), .A3(new_n915), .ZN(new_n923));
  XNOR2_X1  g722(.A(KEYINPUT125), .B(G204gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR4_X1   g724(.A1(new_n837), .A2(new_n651), .A3(new_n918), .A4(new_n924), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1353gat));
  NAND4_X1  g727(.A1(new_n876), .A2(new_n551), .A3(new_n877), .A4(new_n915), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n931), .A2(G211gat), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n362), .A3(new_n551), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n914), .A2(new_n930), .A3(new_n551), .A4(new_n915), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n940), .A3(G211gat), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n934), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n938), .A3(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n916), .B2(new_n731), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n919), .A2(new_n363), .A3(new_n604), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


