//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G15gat), .ZN(new_n204));
  INV_X1    g003(.A(G15gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n206), .C1(new_n207), .C2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(G1gat), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI221_X1 g012(.A(new_n208), .B1(new_n209), .B2(new_n202), .C1(G1gat), .C2(new_n211), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(KEYINPUT14), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT15), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(G43gat), .A2(G50gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT14), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n218), .A2(new_n221), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G29gat), .ZN(new_n231));
  INV_X1    g030(.A(G36gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT14), .ZN(new_n233));
  NAND2_X1  g032(.A1(G29gat), .A2(G36gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n226), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT15), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT89), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n243), .B(KEYINPUT17), .C1(new_n230), .C2(new_n237), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n215), .B(new_n239), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n213), .A2(new_n214), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT18), .B1(new_n249), .B2(KEYINPUT91), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(new_n251), .A3(new_n247), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n245), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n248), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n215), .A2(new_n238), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n247), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n248), .B(KEYINPUT13), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G141gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G169gat), .B(G197gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT12), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n259), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n253), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n250), .B2(new_n252), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(new_n267), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT35), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT84), .B(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277));
  INV_X1    g076(.A(G141gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(G148gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G155gat), .ZN(new_n283));
  INV_X1    g082(.A(G155gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n286), .ZN(new_n288));
  AND2_X1   g087(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n289), .A2(new_n290), .A3(new_n278), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(new_n279), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT77), .B(G162gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n277), .B1(new_n293), .B2(G155gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n287), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT78), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n296));
  OR2_X1    g095(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(G141gat), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n278), .A2(G148gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n286), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(KEYINPUT77), .A2(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(G155gat), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n301), .A2(new_n305), .B1(new_n286), .B2(new_n281), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT29), .B1(new_n296), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(KEYINPUT22), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  NOR2_X1   g116(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n315), .B(new_n316), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n308), .B1(new_n320), .B2(KEYINPUT29), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n321), .B2(new_n295), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT83), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(new_n325), .C1(new_n310), .C2(new_n317), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT3), .B1(new_n317), .B2(new_n332), .ZN(new_n333));
  AOI221_X4 g132(.A(KEYINPUT79), .B1(new_n281), .B2(new_n286), .C1(new_n301), .C2(new_n305), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n301), .A2(new_n305), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n287), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n319), .B1(new_n318), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n327), .A2(new_n331), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n331), .B1(new_n327), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n276), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n330), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n331), .A3(new_n340), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n275), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT23), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT65), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n354), .A2(new_n356), .A3(new_n359), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT66), .B1(new_n349), .B2(KEYINPUT23), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n365), .B(new_n366), .C1(G169gat), .C2(G176gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT68), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n357), .A2(new_n372), .A3(new_n358), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n357), .B2(new_n358), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n353), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT70), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT69), .B(G190gat), .Z(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(G183gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT69), .B(G190gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(KEYINPUT70), .A3(new_n360), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT67), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n350), .A2(new_n382), .A3(new_n351), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n350), .B2(new_n351), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT25), .B(new_n368), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n371), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  OR3_X1    g187(.A1(new_n387), .A2(new_n349), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n387), .B2(new_n349), .ZN(new_n390));
  INV_X1    g189(.A(new_n349), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n389), .B(new_n390), .C1(KEYINPUT26), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n379), .A2(KEYINPUT28), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G183gat), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n394), .A2(new_n396), .A3(KEYINPUT72), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT72), .B1(new_n394), .B2(new_n396), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n394), .A2(new_n396), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n357), .B(new_n392), .C1(new_n399), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n405));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(KEYINPUT1), .ZN(new_n408));
  INV_X1    g207(.A(G120gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G113gat), .ZN(new_n410));
  INV_X1    g209(.A(G113gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G120gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT1), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(G127gat), .A2(G134gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(G127gat), .A2(G134gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n404), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT64), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n408), .A2(new_n417), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n386), .A2(new_n422), .A3(new_n403), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT34), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT75), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n430), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n424), .B(KEYINPUT32), .C1(new_n426), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n431), .B2(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n423), .ZN(new_n440));
  INV_X1    g239(.A(new_n421), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n440), .A2(new_n441), .B1(KEYINPUT75), .B2(new_n432), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n431), .A2(new_n436), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n433), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(new_n437), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n348), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n296), .A2(new_n309), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n418), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n295), .A2(new_n422), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT80), .B1(new_n306), .B2(new_n418), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n295), .A2(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n306), .A2(new_n335), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT4), .A4(new_n418), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n456), .A2(new_n457), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n459), .B1(new_n295), .B2(new_n422), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n306), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n468), .A2(new_n469), .B1(new_n295), .B2(new_n422), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n460), .A2(new_n461), .B1(new_n306), .B2(new_n418), .ZN(new_n472));
  INV_X1    g271(.A(new_n457), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n474));
  AND4_X1   g273(.A1(KEYINPUT5), .A2(new_n466), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n476), .A3(new_n457), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT4), .B1(new_n338), .B2(new_n418), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n460), .A2(new_n461), .A3(new_n458), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n418), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n458), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT4), .A3(new_n469), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(KEYINPUT82), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n477), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n453), .B1(new_n475), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n466), .A2(KEYINPUT5), .A3(new_n471), .A4(new_n474), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n483), .A2(KEYINPUT82), .A3(new_n484), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT82), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n489), .B(new_n452), .C1(new_n492), .C2(new_n477), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT6), .B(new_n453), .C1(new_n475), .C2(new_n486), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G226gat), .ZN(new_n497));
  INV_X1    g296(.A(G233gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n404), .B2(new_n332), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n497), .B(new_n498), .C1(new_n386), .C2(new_n403), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n320), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n404), .A2(new_n499), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n386), .B2(new_n403), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n503), .B(new_n317), .C1(new_n499), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n507), .B(new_n508), .Z(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n502), .A2(new_n509), .A3(new_n505), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n512), .ZN(new_n513));
  OR3_X1    g312(.A1(new_n506), .A2(KEYINPUT30), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n274), .B1(new_n448), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n443), .B1(new_n438), .B2(new_n439), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n446), .A2(new_n442), .A3(new_n437), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n518), .A2(new_n519), .B1(new_n343), .B2(new_n347), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n494), .A2(new_n495), .B1(new_n514), .B2(new_n513), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(KEYINPUT87), .A3(KEYINPUT35), .A4(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT36), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT36), .B1(new_n518), .B2(new_n519), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n348), .ZN(new_n528));
  INV_X1    g327(.A(new_n496), .ZN(new_n529));
  INV_X1    g328(.A(new_n515), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT39), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n470), .B2(new_n457), .ZN(new_n533));
  INV_X1    g332(.A(new_n456), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n481), .B2(new_n485), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(new_n457), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n456), .B1(new_n490), .B2(new_n491), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n532), .A3(new_n473), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n452), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n539), .A2(KEYINPUT85), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n539), .B2(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n487), .A2(new_n513), .A3(new_n514), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n502), .A2(new_n545), .A3(new_n505), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT37), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n502), .A2(new_n545), .A3(new_n505), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n510), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT38), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT38), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n547), .A2(new_n552), .A3(new_n510), .A4(new_n549), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n512), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n348), .B1(new_n554), .B2(new_n496), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n527), .B(new_n531), .C1(new_n544), .C2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n273), .B1(new_n523), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G57gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G64gat), .ZN(new_n565));
  INV_X1    g364(.A(G64gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(G57gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G127gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n215), .B1(new_n573), .B2(new_n572), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT93), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n582), .B(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n590), .A2(new_n593), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n240), .B2(new_n241), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n243), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n240), .A2(KEYINPUT89), .A3(new_n241), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n598), .A2(new_n600), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n614), .A2(new_n240), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(G190gat), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n242), .A2(new_n244), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n361), .B(new_n617), .C1(new_n620), .C2(new_n608), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT95), .B1(new_n622), .B2(new_n313), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(G218gat), .A3(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT94), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n588), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n572), .B1(new_n612), .B2(new_n613), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n601), .A2(new_n563), .A3(new_n606), .A4(new_n571), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n563), .A4(new_n571), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n635), .A2(new_n637), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G120gat), .B(G148gat), .Z(new_n647));
  XOR2_X1   g446(.A(G176gat), .B(G204gat), .Z(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(new_n645), .A3(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n634), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n557), .A2(new_n529), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT96), .B(G1gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n557), .A2(new_n656), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n530), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT42), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n660), .B2(new_n515), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT97), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(KEYINPUT97), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n660), .B2(new_n527), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n444), .A2(new_n447), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n205), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n669), .B1(new_n660), .B2(new_n672), .ZN(G1326gat));
  OR3_X1    g472(.A1(new_n660), .A2(KEYINPUT98), .A3(new_n348), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT98), .B1(new_n660), .B2(new_n348), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(new_n588), .ZN(new_n679));
  INV_X1    g478(.A(new_n633), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n679), .A2(new_n680), .A3(new_n653), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n557), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n496), .A2(G29gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT99), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n686), .A2(KEYINPUT45), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT45), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n544), .A2(new_n555), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT36), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n444), .B2(new_n447), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n524), .C1(new_n348), .C2(new_n521), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n517), .B(new_n522), .C1(new_n693), .C2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n633), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n697), .B2(new_n633), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n588), .B(KEYINPUT100), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n273), .A3(new_n653), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n692), .B1(new_n704), .B2(new_n496), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n701), .A2(KEYINPUT101), .A3(new_n529), .A4(new_n703), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(G29gat), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n707), .ZN(G1328gat));
  NOR3_X1   g507(.A1(new_n682), .A2(G36gat), .A3(new_n515), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n704), .B2(new_n515), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  NAND3_X1  g511(.A1(new_n557), .A2(new_n671), .A3(new_n681), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n713), .A2(new_n222), .B1(KEYINPUT102), .B2(KEYINPUT47), .ZN(new_n714));
  INV_X1    g513(.A(new_n527), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n704), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1330gat));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n633), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n722), .A2(new_n528), .A3(new_n698), .A4(new_n703), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n683), .A2(new_n223), .A3(new_n528), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1331gat));
  NAND3_X1  g527(.A1(new_n634), .A2(new_n273), .A3(new_n653), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n523), .B2(new_n556), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n529), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g531(.A(new_n515), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT103), .Z(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n730), .A2(new_n738), .A3(new_n671), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n730), .A2(new_n715), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n738), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g541(.A1(new_n730), .A2(new_n528), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT104), .B(G78gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  XNOR2_X1  g544(.A(new_n271), .B(new_n267), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n679), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n653), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT105), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n701), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n496), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n693), .A2(new_n696), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n517), .A2(new_n522), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n633), .B(new_n747), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n697), .A2(KEYINPUT51), .A3(new_n633), .A4(new_n747), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n529), .A2(new_n594), .A3(new_n653), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n751), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NAND2_X1  g560(.A1(new_n530), .A2(new_n653), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n680), .B1(new_n523), .B2(new_n556), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT51), .B1(new_n764), .B2(new_n747), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n722), .A2(new_n530), .A3(new_n698), .A4(new_n749), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n758), .A2(KEYINPUT107), .A3(new_n763), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n776), .B(new_n777), .C1(new_n767), .C2(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1337gat));
  NOR2_X1   g578(.A1(new_n750), .A2(new_n527), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT108), .B(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n671), .A2(new_n653), .A3(new_n781), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n780), .A2(new_n781), .B1(new_n759), .B2(new_n782), .ZN(G1338gat));
  NAND4_X1  g582(.A1(new_n722), .A2(new_n528), .A3(new_n698), .A4(new_n749), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n348), .A2(G106gat), .A3(new_n654), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT109), .B1(new_n758), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  INV_X1    g587(.A(new_n786), .ZN(new_n789));
  AOI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n756), .C2(new_n757), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n785), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT53), .B1(new_n758), .B2(new_n786), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n784), .A2(G106gat), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n793), .A2(KEYINPUT110), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT110), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n792), .B1(new_n795), .B2(new_n796), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n656), .A2(new_n273), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  INV_X1    g598(.A(new_n266), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n245), .A2(new_n247), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n801), .A2(new_n248), .B1(new_n257), .B2(new_n258), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n271), .A2(new_n800), .B1(new_n265), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n629), .B1(new_n623), .B2(new_n624), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n807));
  AND4_X1   g606(.A1(KEYINPUT111), .A2(new_n642), .A3(KEYINPUT54), .A4(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n640), .B2(new_n641), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT111), .B1(new_n810), .B2(new_n807), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n644), .B1(new_n638), .B2(new_n639), .ZN(new_n813));
  AOI211_X1 g612(.A(new_n812), .B(new_n649), .C1(new_n813), .C2(new_n809), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n640), .A2(new_n809), .A3(new_n641), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n815), .B2(new_n650), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n808), .A2(new_n811), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI211_X1 g618(.A(KEYINPUT54), .B(new_n644), .C1(new_n638), .C2(new_n639), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n812), .B1(new_n820), .B2(new_n649), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(KEYINPUT112), .A3(new_n650), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(KEYINPUT55), .C1(new_n811), .C2(new_n808), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n819), .A2(new_n652), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n799), .B1(new_n806), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n819), .A2(new_n652), .A3(new_n824), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(new_n633), .A3(KEYINPUT113), .A4(new_n803), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n803), .A2(new_n653), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n830), .B(new_n831), .C1(new_n273), .C2(new_n825), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n273), .B2(new_n825), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n633), .B1(new_n833), .B2(KEYINPUT114), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n829), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n798), .B1(new_n835), .B2(new_n702), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n348), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n496), .A2(new_n530), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n671), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n273), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n836), .A2(new_n529), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n520), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n530), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT115), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n746), .A2(new_n411), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n839), .B2(new_n654), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n653), .A2(new_n409), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n844), .B2(new_n849), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n577), .A3(new_n679), .ZN(new_n851));
  INV_X1    g650(.A(new_n702), .ZN(new_n852));
  OAI21_X1  g651(.A(G127gat), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1342gat));
  NAND2_X1  g653(.A1(new_n633), .A2(new_n515), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT117), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n842), .A2(G134gat), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n839), .B2(new_n680), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n715), .A2(new_n348), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n530), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n273), .A2(G141gat), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT120), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n527), .A2(new_n838), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n836), .B2(new_n528), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n528), .A2(KEYINPUT57), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n826), .A2(new_n828), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n253), .A2(new_n269), .A3(new_n800), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n802), .A2(new_n265), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n875), .A2(new_n653), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n827), .B2(new_n746), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n680), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n833), .A2(KEYINPUT119), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n588), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n873), .B1(new_n883), .B2(new_n798), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n869), .B1(new_n872), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT121), .B1(new_n885), .B2(new_n273), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n273), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n867), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n864), .A2(new_n866), .ZN(new_n890));
  INV_X1    g689(.A(new_n885), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n278), .B1(new_n891), .B2(new_n746), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT58), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n289), .A2(new_n290), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n864), .A2(new_n895), .A3(new_n653), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n895), .C1(new_n891), .C2(new_n653), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n655), .A2(new_n746), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n806), .A2(new_n825), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n880), .B2(new_n881), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(new_n588), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n899), .B1(new_n904), .B2(new_n348), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n833), .A2(KEYINPUT114), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n680), .A3(new_n832), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n702), .B1(new_n907), .B2(new_n874), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n528), .B(new_n871), .C1(new_n908), .C2(new_n900), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n653), .A3(new_n869), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n898), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n864), .A2(new_n284), .A3(new_n679), .ZN(new_n914));
  OAI21_X1  g713(.A(G155gat), .B1(new_n885), .B2(new_n852), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(new_n293), .B1(new_n885), .B2(new_n680), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n856), .A2(new_n293), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n863), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n529), .A2(new_n515), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n670), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n837), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(G169gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n273), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n836), .A2(new_n496), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n448), .A2(new_n515), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n746), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n924), .B2(new_n930), .ZN(G1348gat));
  INV_X1    g730(.A(G176gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n923), .A2(new_n932), .A3(new_n654), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n653), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(G1349gat));
  OAI21_X1  g734(.A(G183gat), .B1(new_n923), .B2(new_n852), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n588), .A2(new_n398), .A3(new_n397), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(G1350gat));
  NOR3_X1   g739(.A1(new_n928), .A2(new_n377), .A3(new_n680), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n837), .A2(new_n633), .A3(new_n922), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT123), .B1(new_n943), .B2(G190gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(new_n942), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n943), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n910), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n905), .A2(KEYINPUT124), .A3(new_n909), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n715), .A2(new_n921), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n273), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n926), .A2(new_n862), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n746), .A3(new_n530), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n954), .A2(new_n956), .B1(new_n959), .B2(new_n955), .ZN(G1352gat));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  AOI211_X1 g760(.A(G204gat), .B(new_n762), .C1(new_n961), .C2(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n963), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(G204gat), .B1(new_n953), .B2(new_n654), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1353gat));
  NAND4_X1  g766(.A1(new_n958), .A2(new_n312), .A3(new_n530), .A4(new_n679), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n679), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n905), .B2(new_n909), .ZN(new_n970));
  NAND2_X1  g769(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n971));
  OAI21_X1  g770(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n971), .ZN(new_n974));
  INV_X1    g773(.A(new_n969), .ZN(new_n975));
  INV_X1    g774(.A(new_n909), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n633), .B1(new_n833), .B2(KEYINPUT119), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n878), .A2(new_n879), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n901), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n798), .B1(new_n979), .B2(new_n679), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT57), .B1(new_n980), .B2(new_n528), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n975), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n972), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n968), .B1(new_n973), .B2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g786(.A(KEYINPUT127), .B(new_n968), .C1(new_n973), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1354gat));
  NOR2_X1   g788(.A1(new_n680), .A2(new_n313), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n958), .A2(new_n530), .A3(new_n633), .ZN(new_n991));
  AOI22_X1  g790(.A1(new_n954), .A2(new_n990), .B1(new_n991), .B2(new_n313), .ZN(G1355gat));
endmodule


