//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(new_n457), .B1(G567), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(new_n457), .B2(new_n456), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n459), .B(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n479), .A2(new_n484), .ZN(G162));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(KEYINPUT70), .B2(G114), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT70), .A2(G114), .ZN(new_n488));
  OAI211_X1 g063(.A(G2104), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n463), .B2(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n464), .C2(new_n463), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n504), .B2(KEYINPUT71), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT71), .A3(G62), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n506), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G88), .B1(new_n516), .B2(G50), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n513), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n502), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(new_n516), .A2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(new_n521), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n502), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(new_n539), .B2(new_n538), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT75), .B(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n530), .A2(new_n544), .B1(new_n522), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n535), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n558));
  NAND3_X1  g133(.A1(new_n516), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n514), .A2(G91), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n535), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n502), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n568), .A2(KEYINPUT77), .A3(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n562), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n500), .A2(new_n501), .A3(G74), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n535), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT78), .B(G651), .C1(new_n508), .C2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n514), .A2(G87), .B1(new_n516), .B2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  INV_X1    g156(.A(G73), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n502), .A2(new_n581), .B1(new_n582), .B2(new_n515), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(new_n513), .ZN(new_n585));
  NOR2_X1   g160(.A1(KEYINPUT6), .A2(G651), .ZN(new_n586));
  OAI211_X1 g161(.A(G48), .B(G543), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n583), .A2(G651), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n514), .A2(G86), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n516), .A2(KEYINPUT79), .A3(G48), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n535), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n516), .A2(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n530), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n593), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n514), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT82), .B(G66), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n508), .A2(new_n602), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n535), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G54), .B1(new_n516), .B2(KEYINPUT81), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT83), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n604), .B(new_n610), .C1(new_n606), .C2(new_n607), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n601), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G286), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(G299), .B(KEYINPUT84), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G297));
  AOI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(new_n615), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT85), .ZN(G148));
  NAND2_X1  g197(.A1(new_n612), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g201(.A(KEYINPUT3), .B(G2104), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n470), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  AOI22_X1  g208(.A1(G123), .A2(new_n477), .B1(new_n483), .B2(G135), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n635), .A2(new_n462), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n462), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n643), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g235(.A(KEYINPUT88), .B(new_n658), .C1(new_n655), .C2(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n657), .B2(new_n659), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n631), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n640), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT91), .ZN(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n693), .A2(new_n694), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  AOI22_X1  g281(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n477), .A2(G129), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(G32), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT27), .B(G1996), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT103), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n716), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G116), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G128), .B2(new_n477), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n483), .A2(new_n729), .A3(G140), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n483), .B2(G140), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n724), .B1(new_n733), .B2(new_n716), .ZN(new_n734));
  INV_X1    g309(.A(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G27), .A2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G164), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT104), .B(G2078), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n736), .B(new_n742), .C1(new_n718), .C2(new_n720), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n722), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n716), .A2(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n716), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT29), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G2090), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G19), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n549), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G16), .ZN(new_n754));
  NOR2_X1   g329(.A1(G168), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NAND2_X1  g332(.A1(G160), .A2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n759), .B2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT24), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n756), .A2(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT25), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G139), .B2(new_n483), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n462), .B2(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G33), .B(new_n769), .S(G29), .Z(new_n770));
  AOI211_X1 g345(.A(new_n753), .B(new_n764), .C1(G2072), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G11), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n716), .B1(new_n773), .B2(G28), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n772), .B1(new_n774), .B2(new_n775), .C1(new_n639), .C2(new_n716), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n762), .B2(new_n763), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n756), .A2(new_n757), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G2072), .B2(new_n770), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n752), .B2(new_n751), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n771), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n754), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n754), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1961), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n748), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n754), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G299), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n754), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n747), .B2(G2090), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT106), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n754), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n612), .B2(new_n754), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1348), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n792), .B2(KEYINPUT106), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n744), .A2(new_n786), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n754), .A2(G23), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n578), .A2(new_n579), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n754), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT98), .Z(new_n802));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G1976), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n802), .B(KEYINPUT33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G1976), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n754), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n754), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1971), .ZN(new_n811));
  MUX2_X1   g386(.A(G6), .B(G305), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n806), .A2(new_n808), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  OAI21_X1  g393(.A(KEYINPUT93), .B1(G95), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(KEYINPUT93), .A2(G95), .A3(G2105), .ZN(new_n821));
  OAI221_X1 g396(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(G119), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n627), .A2(G2105), .ZN(new_n824));
  INV_X1    g399(.A(G131), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n627), .A2(new_n462), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT94), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G29), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n716), .A2(G25), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n818), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  INV_X1    g411(.A(new_n818), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n754), .B1(G290), .B2(KEYINPUT96), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(KEYINPUT96), .B2(G290), .ZN(new_n841));
  INV_X1    g416(.A(G24), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(G16), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G1986), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT34), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n806), .A2(new_n808), .A3(new_n851), .A4(new_n815), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n849), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n817), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT36), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(new_n817), .C1(new_n853), .C2(new_n854), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n798), .B1(new_n856), .B2(new_n858), .ZN(G311));
  INV_X1    g434(.A(new_n798), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n849), .A2(new_n852), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n857), .B1(new_n864), .B2(new_n817), .ZN(new_n865));
  INV_X1    g440(.A(new_n858), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(G150));
  NAND2_X1  g442(.A1(new_n612), .A2(G559), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT38), .Z(new_n869));
  AOI22_X1  g444(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n535), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n516), .A2(G55), .ZN(new_n872));
  INV_X1    g447(.A(G93), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n530), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n548), .B2(new_n546), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n871), .A2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n549), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n869), .B(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n877), .A2(new_n882), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(G145));
  NAND2_X1  g462(.A1(new_n495), .A2(new_n497), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT70), .ZN(new_n889));
  INV_X1    g464(.A(G114), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(KEYINPUT70), .A2(G114), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(G2105), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(G126), .A2(new_n477), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n714), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n714), .A2(new_n897), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n827), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n769), .A2(new_n732), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n483), .A2(G142), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n477), .A2(G130), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n462), .A2(G118), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n629), .B(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n769), .A2(new_n732), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n903), .B2(new_n910), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n899), .A2(new_n827), .A3(new_n900), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n902), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  INV_X1    g491(.A(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n901), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n639), .B(G160), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G162), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n915), .A2(new_n918), .A3(new_n921), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g502(.A1(new_n875), .A2(new_n615), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n609), .A2(new_n611), .ZN(new_n929));
  INV_X1    g504(.A(new_n601), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n612), .A2(new_n789), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT41), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n623), .B(new_n879), .Z(new_n939));
  MUX2_X1   g514(.A(new_n935), .B(new_n938), .S(new_n939), .Z(new_n940));
  NOR2_X1   g515(.A1(new_n593), .A2(new_n596), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT107), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(G288), .ZN(new_n943));
  XNOR2_X1  g518(.A(G166), .B(G305), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n940), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n928), .B1(new_n947), .B2(new_n615), .ZN(G295));
  OAI21_X1  g523(.A(new_n928), .B1(new_n947), .B2(new_n615), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n934), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n952));
  NAND2_X1  g527(.A1(G171), .A2(new_n879), .ZN(new_n953));
  NAND3_X1  g528(.A1(G301), .A2(new_n876), .A3(new_n878), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(G168), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n954), .ZN(new_n956));
  AOI21_X1  g531(.A(G301), .B1(new_n876), .B2(new_n878), .ZN(new_n957));
  OAI21_X1  g532(.A(G286), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n951), .A2(new_n952), .A3(new_n955), .A4(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n955), .ZN(new_n960));
  AOI21_X1  g535(.A(G168), .B1(new_n953), .B2(new_n954), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n935), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n945), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n924), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n960), .A2(new_n961), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n938), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n962), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n934), .B1(new_n958), .B2(new_n955), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n966), .A2(new_n969), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n972), .B1(new_n938), .B2(new_n967), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n945), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n963), .A2(new_n964), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT43), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n978), .B2(new_n979), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n975), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(KEYINPUT44), .B2(new_n984), .ZN(G397));
  INV_X1    g560(.A(KEYINPUT126), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  INV_X1    g562(.A(new_n497), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n496), .B1(new_n627), .B2(new_n493), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n987), .B1(new_n990), .B2(new_n491), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  INV_X1    g567(.A(G40), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n467), .A2(new_n472), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n715), .B2(G1996), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n714), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n827), .B(KEYINPUT112), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n995), .B1(new_n1000), .B2(new_n837), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n837), .B2(new_n1000), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n732), .A2(G2067), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n732), .A2(G2067), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1006), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT110), .A3(new_n1004), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n995), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT111), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1013), .B(new_n995), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n999), .B(new_n1002), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n941), .A2(new_n846), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n995), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  NAND2_X1  g595(.A1(G160), .A2(G40), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n888), .B2(new_n896), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1023), .A2(new_n1026), .A3(new_n1022), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1024), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1961), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1021), .B1(new_n991), .B2(new_n992), .ZN(new_n1031));
  INV_X1    g606(.A(G2078), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n897), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(KEYINPUT53), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1035), .A2(new_n1032), .A3(new_n1033), .A4(new_n994), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1030), .A2(G301), .A3(new_n1034), .A4(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1022), .B(new_n987), .C1(new_n990), .C2(new_n491), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n994), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1026), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n991), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1038), .B(new_n1034), .C1(new_n1044), .C2(G1961), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(G171), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1045), .B2(G171), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1039), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n994), .B1(new_n1023), .B2(KEYINPUT45), .ZN(new_n1052));
  NOR3_X1   g627(.A1(G164), .A2(new_n992), .A3(G1384), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n757), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n763), .B(new_n1024), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT119), .B(new_n757), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(G286), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(G168), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1061), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1045), .A2(G171), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT54), .A3(new_n1039), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1023), .A2(new_n994), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n578), .A2(new_n1071), .A3(G1976), .A4(new_n579), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1070), .A2(G8), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT115), .B1(G288), .B2(new_n805), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1976), .B1(new_n578), .B2(new_n579), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT116), .B1(new_n1075), .B2(KEYINPUT52), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(new_n1078), .C1(new_n800), .C2(G1976), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1981), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n588), .A2(new_n1081), .A3(new_n589), .A4(new_n590), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT117), .B(G86), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n514), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n581), .B1(new_n506), .B2(new_n507), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n582), .A2(new_n515), .ZN(new_n1086));
  OAI21_X1  g661(.A(G651), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n587), .A2(new_n584), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n590), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1023), .B2(new_n994), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1082), .A2(new_n1090), .A3(KEYINPUT49), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1072), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1074), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1080), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G166), .A2(new_n1094), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT55), .ZN(new_n1103));
  INV_X1    g678(.A(G2090), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1024), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1105));
  INV_X1    g680(.A(G1971), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1094), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(new_n1104), .A3(new_n994), .A4(new_n1040), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1111), .A3(KEYINPUT118), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(G8), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1102), .B(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1069), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1051), .A2(new_n1067), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1051), .A2(new_n1067), .A3(new_n1120), .A4(KEYINPUT122), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1070), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n1023), .B2(new_n994), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1128), .A2(new_n735), .B1(new_n1028), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT58), .B(G1341), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1126), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1052), .A2(new_n1053), .A3(G1996), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n549), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT59), .B(new_n549), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n562), .A2(new_n570), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n562), .B2(new_n570), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1956), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1023), .A2(new_n1022), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1041), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1031), .A2(new_n1033), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1144), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1144), .A2(new_n1149), .A3(new_n1147), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT61), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1152), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1154), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1140), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1130), .B(new_n931), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT60), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1130), .A2(new_n931), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1150), .B1(new_n1161), .B2(new_n1152), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1123), .A2(new_n1124), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1059), .A2(G286), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1065), .B1(new_n1064), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1063), .A2(new_n1066), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1048), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1045), .A2(new_n1046), .A3(G171), .ZN(new_n1172));
  AND4_X1   g747(.A1(new_n1171), .A2(new_n1109), .A3(new_n1119), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1095), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1082), .ZN(new_n1177));
  NOR2_X1   g752(.A1(G288), .A2(G1976), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1097), .B2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1175), .A2(new_n1101), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1059), .A2(G8), .A3(G168), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1109), .A2(new_n1119), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1185), .A2(new_n1109), .A3(KEYINPUT63), .A4(new_n1181), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1180), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1020), .B1(new_n1164), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n828), .A2(new_n837), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n999), .B(new_n1190), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1008), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT123), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1191), .A2(new_n1194), .A3(new_n1008), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1193), .A2(new_n1011), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1193), .A2(KEYINPUT124), .A3(new_n1011), .A4(new_n1195), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1011), .A2(new_n997), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT46), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1011), .B1(new_n1010), .B2(new_n714), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT47), .Z(new_n1205));
  NOR2_X1   g780(.A1(new_n995), .A2(new_n1017), .ZN(new_n1206));
  XOR2_X1   g781(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1207));
  NOR2_X1   g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AND2_X1   g783(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1015), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1205), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1200), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n986), .B1(new_n1189), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1211), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1216));
  AOI22_X1  g791(.A1(new_n1121), .A2(new_n1122), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n1217), .B2(new_n1124), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1215), .B(KEYINPUT126), .C1(new_n1218), .C2(new_n1020), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1213), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n1222));
  INV_X1    g796(.A(G227), .ZN(new_n1223));
  NAND2_X1  g797(.A1(G319), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1224), .B1(new_n662), .B2(new_n664), .ZN(new_n1225));
  NAND3_X1  g799(.A1(new_n705), .A2(new_n926), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n974), .A2(new_n964), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n1227), .A2(new_n982), .A3(new_n978), .ZN(new_n1228));
  NAND2_X1  g802(.A1(new_n978), .A2(new_n979), .ZN(new_n1229));
  NAND2_X1  g803(.A1(new_n1229), .A2(KEYINPUT43), .ZN(new_n1230));
  AOI211_X1 g804(.A(new_n1222), .B(new_n1226), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1232));
  INV_X1    g806(.A(new_n1226), .ZN(new_n1233));
  AOI21_X1  g807(.A(KEYINPUT127), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n1231), .A2(new_n1234), .ZN(G308));
  OAI21_X1  g809(.A(new_n1222), .B1(new_n984), .B2(new_n1226), .ZN(new_n1236));
  NAND3_X1  g810(.A1(new_n1232), .A2(KEYINPUT127), .A3(new_n1233), .ZN(new_n1237));
  NAND2_X1  g811(.A1(new_n1236), .A2(new_n1237), .ZN(G225));
endmodule


