//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1192, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT64), .Z(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n225), .A2(new_n226), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  AOI21_X1  g0051(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT66), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(G222), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n217), .B2(new_n257), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n252), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT65), .B1(new_n253), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n230), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G33), .A3(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G274), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(G226), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n265), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT67), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n265), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G190), .ZN(new_n285));
  XOR2_X1   g0085(.A(KEYINPUT8), .B(G58), .Z(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n288), .B1(G150), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(G20), .B2(new_n203), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n291), .B2(new_n290), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n230), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n207), .A3(G1), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n206), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G50), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n296), .B(new_n301), .C1(G50), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT9), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n281), .A2(new_n283), .A3(G200), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n285), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n285), .A2(new_n304), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n284), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n303), .C1(G169), .C2(new_n284), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G77), .B2(new_n302), .ZN(new_n316));
  INV_X1    g0116(.A(new_n295), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n286), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n288), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n259), .A2(new_n212), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n257), .A2(G232), .A3(new_n262), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n254), .A2(new_n256), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT71), .B(G107), .Z(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n326), .B2(new_n325), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n252), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n274), .B1(new_n277), .B2(new_n218), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G179), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n323), .B1(new_n338), .B2(KEYINPUT72), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n340), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n339), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(G190), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n323), .C1(new_n345), .C2(new_n337), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n237), .A2(G1698), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G226), .B2(G1698), .ZN(new_n349));
  INV_X1    g0149(.A(G97), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n327), .B1(new_n253), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n252), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n274), .C1(new_n212), .C2(new_n277), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT13), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n298), .A2(new_n211), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n217), .B2(new_n287), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT11), .B1(new_n361), .B2(new_n295), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n354), .B2(new_n345), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n354), .A2(G169), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n355), .A2(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n366), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n314), .A2(new_n347), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n255), .B2(G33), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n253), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n256), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n260), .A2(new_n262), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G226), .B2(new_n262), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n383), .A2(new_n385), .B1(new_n253), .B2(new_n213), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI221_X1 g0188(.A(KEYINPUT78), .B1(new_n253), .B2(new_n213), .C1(new_n383), .C2(new_n385), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n252), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n277), .A2(new_n237), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(new_n275), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n341), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n390), .A2(new_n392), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(G179), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n383), .A2(new_n207), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n211), .B1(new_n398), .B2(KEYINPUT7), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n383), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n381), .A2(new_n382), .A3(KEYINPUT75), .A4(new_n256), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT7), .A2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT76), .B1(new_n399), .B2(new_n404), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n397), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n327), .A2(new_n207), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT7), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n397), .B1(new_n409), .B2(new_n211), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n407), .A2(new_n412), .A3(new_n295), .ZN(new_n413));
  INV_X1    g0213(.A(new_n299), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n286), .A2(new_n300), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n414), .A2(new_n415), .B1(new_n302), .B2(new_n286), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n395), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n356), .B1(new_n390), .B2(new_n392), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(G190), .B2(new_n394), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n413), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT79), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n413), .A2(new_n422), .A3(new_n417), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(new_n425), .A3(new_n426), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n420), .A2(new_n428), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n379), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n271), .A2(G274), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n272), .A2(G1), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  NOR2_X1   g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n271), .A2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G264), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n214), .A2(new_n262), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G257), .B2(new_n262), .ZN(new_n446));
  INV_X1    g0246(.A(G294), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n383), .A2(new_n446), .B1(new_n253), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n252), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n442), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G190), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n449), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT84), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n455), .B2(new_n356), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT23), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n219), .A3(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n458), .B1(KEYINPUT83), .B2(new_n459), .C1(new_n460), .C2(new_n287), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n257), .A2(new_n207), .A3(G87), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT23), .B1(new_n329), .B2(new_n207), .ZN(new_n465));
  INV_X1    g0265(.A(new_n383), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n207), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT22), .A2(G87), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n464), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n295), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n297), .A2(G1), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G20), .A3(new_n219), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT25), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n299), .B1(G1), .B2(new_n253), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(G107), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n456), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n450), .A2(G169), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n455), .B2(new_n311), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n479), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT7), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n408), .B(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT6), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n350), .A2(new_n219), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n486), .A2(new_n329), .B1(new_n493), .B2(KEYINPUT80), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n493), .A2(KEYINPUT80), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n295), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n298), .A2(new_n350), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n476), .B2(new_n350), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n443), .A2(G257), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n442), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n214), .B2(new_n262), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n257), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n383), .A2(new_n218), .A3(G1698), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n506), .B(new_n509), .C1(new_n510), .C2(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n252), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n442), .A2(new_n502), .A3(KEYINPUT81), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n505), .A2(new_n311), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n505), .A2(new_n513), .A3(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n341), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n501), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n499), .B1(new_n496), .B2(new_n295), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(G200), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n345), .C2(new_n515), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n443), .A2(G270), .ZN(new_n522));
  INV_X1    g0322(.A(new_n252), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G257), .A2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n220), .B2(G1698), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n466), .A2(new_n525), .B1(G303), .B2(new_n327), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n442), .B(new_n522), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n506), .B(new_n207), .C1(G33), .C2(new_n350), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(new_n295), .C1(new_n207), .C2(G116), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n298), .A2(new_n460), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n476), .B2(new_n460), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OR3_X1    g0334(.A1(new_n528), .A2(KEYINPUT21), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT21), .B1(new_n528), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n534), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G200), .B2(new_n527), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n345), .B2(new_n527), .ZN(new_n540));
  INV_X1    g0340(.A(new_n527), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n538), .A2(new_n541), .A3(G179), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n328), .A2(new_n213), .A3(new_n350), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n207), .B1(new_n253), .B2(new_n350), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n287), .A2(KEYINPUT19), .A3(new_n350), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(new_n211), .B2(new_n467), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(new_n295), .B1(new_n298), .B2(new_n319), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n477), .A2(new_n320), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OR3_X1    g0352(.A1(new_n272), .A2(G1), .A3(G274), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n271), .B(new_n553), .C1(G250), .C2(new_n438), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT82), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n218), .A2(G1698), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G238), .B2(G1698), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n383), .A2(new_n557), .B1(new_n253), .B2(new_n460), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n252), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n311), .ZN(new_n561));
  INV_X1    g0361(.A(new_n559), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(KEYINPUT82), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n341), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n552), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n356), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n477), .A2(G87), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n550), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n543), .A2(new_n572), .ZN(new_n573));
  AND4_X1   g0373(.A1(new_n436), .A2(new_n484), .A3(new_n521), .A4(new_n573), .ZN(G372));
  OAI21_X1  g0374(.A(new_n377), .B1(new_n343), .B2(new_n368), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n575), .A2(new_n428), .A3(new_n432), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n420), .A2(new_n430), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n310), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n313), .ZN(new_n579));
  INV_X1    g0379(.A(new_n552), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n561), .B2(new_n566), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n565), .A2(G179), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(KEYINPUT85), .C1(new_n341), .C2(new_n565), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n560), .A2(KEYINPUT86), .A3(G200), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n565), .B2(new_n356), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(new_n571), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n585), .A2(new_n517), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT88), .B1(new_n591), .B2(KEYINPUT26), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n582), .A2(new_n584), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n552), .ZN(new_n594));
  INV_X1    g0394(.A(new_n517), .ZN(new_n595));
  INV_X1    g0395(.A(new_n590), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n572), .A2(new_n517), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT26), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n592), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n517), .B(new_n520), .C1(new_n456), .C2(new_n479), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n604), .A2(new_n585), .A3(new_n590), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT87), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n537), .A2(new_n606), .A3(new_n542), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n537), .B2(new_n542), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n483), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n585), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n579), .B1(new_n435), .B2(new_n612), .ZN(G369));
  NAND2_X1  g0413(.A1(new_n473), .A2(new_n207), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(KEYINPUT27), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(KEYINPUT27), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(G213), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g0417(.A(KEYINPUT89), .B(G343), .Z(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n534), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OR3_X1    g0422(.A1(new_n607), .A2(new_n608), .A3(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n537), .A2(new_n542), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n540), .A3(new_n622), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(KEYINPUT90), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n623), .B2(new_n625), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n479), .A2(new_n619), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n484), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n483), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n619), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n632), .A2(G330), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n620), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n624), .A2(new_n619), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n484), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(G399));
  NOR2_X1   g0442(.A1(new_n545), .A2(G116), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n227), .A2(new_n266), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G1), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n233), .B2(new_n644), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT28), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n597), .A2(KEYINPUT26), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n585), .B1(new_n601), .B2(new_n599), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n585), .A2(new_n590), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n480), .A3(new_n521), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n624), .A2(new_n483), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n619), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT29), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n648), .B(new_n649), .C1(new_n652), .C2(new_n653), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n620), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT29), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT91), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n619), .B1(new_n603), .B2(new_n610), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n657), .B(new_n661), .C1(new_n662), .C2(KEYINPUT29), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n484), .A2(new_n521), .A3(new_n573), .A4(new_n620), .ZN(new_n664));
  INV_X1    g0464(.A(new_n515), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(new_n561), .A3(new_n454), .A4(new_n541), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT30), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n541), .A2(new_n565), .A3(G179), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n455), .A2(new_n669), .A3(new_n515), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n619), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT31), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(KEYINPUT31), .A3(new_n619), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n664), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n663), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n647), .B1(new_n680), .B2(G1), .ZN(G364));
  NOR2_X1   g0481(.A1(G13), .A2(G33), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G20), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT93), .Z(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n623), .A2(new_n625), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n230), .B1(G20), .B2(new_n341), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n233), .A2(G45), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n401), .A2(new_n402), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n227), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n690), .B(new_n693), .C1(G45), .C2(new_n250), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n227), .A2(new_n257), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(KEYINPUT92), .B2(G355), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(KEYINPUT92), .B2(G355), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G116), .B2(new_n227), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n689), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n297), .A2(G20), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n206), .B1(new_n700), .B2(G45), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n644), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n207), .A2(new_n311), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G190), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G311), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n207), .A2(G179), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n704), .ZN(new_n708));
  INV_X1    g0508(.A(G329), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n705), .A2(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(G190), .A3(new_n356), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n257), .B(new_n710), .C1(G322), .C2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n345), .A2(G179), .A3(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n207), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n703), .A2(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n345), .ZN(new_n718));
  AOI22_X1  g0518(.A1(G294), .A2(new_n716), .B1(new_n718), .B2(G326), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(G190), .ZN(new_n720));
  XNOR2_X1  g0520(.A(KEYINPUT33), .B(G317), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n707), .A2(new_n345), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n720), .A2(new_n721), .B1(new_n723), .B2(G283), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n713), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n707), .A2(G190), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G303), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n708), .ZN(new_n733));
  XNOR2_X1  g0533(.A(KEYINPUT94), .B(G159), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT95), .B(KEYINPUT32), .Z(new_n736));
  XNOR2_X1  g0536(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n716), .A2(G97), .B1(new_n723), .B2(G107), .ZN(new_n738));
  AOI22_X1  g0538(.A1(G50), .A2(new_n718), .B1(new_n720), .B2(G68), .ZN(new_n739));
  INV_X1    g0539(.A(G58), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n257), .B1(new_n711), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n705), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(G77), .B2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n730), .A2(new_n213), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n725), .A2(new_n732), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n702), .B1(new_n746), .B2(new_n688), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n687), .A2(new_n699), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n627), .B2(new_n630), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n702), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n628), .A2(new_n753), .A3(new_n631), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n748), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(G396));
  NOR2_X1   g0556(.A1(new_n620), .A2(new_n323), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n339), .B(new_n757), .C1(new_n338), .C2(new_n342), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n347), .B2(new_n757), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n662), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n751), .B1(new_n760), .B2(new_n678), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n678), .B2(new_n760), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n711), .A2(new_n447), .B1(new_n708), .B2(new_n706), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n257), .B(new_n763), .C1(G116), .C2(new_n742), .ZN(new_n764));
  INV_X1    g0564(.A(new_n730), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G107), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G97), .A2(new_n716), .B1(new_n718), .B2(G303), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n720), .A2(G283), .B1(new_n723), .B2(G87), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n764), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n712), .A2(G143), .B1(new_n742), .B2(new_n734), .ZN(new_n770));
  INV_X1    g0570(.A(new_n718), .ZN(new_n771));
  INV_X1    g0571(.A(G137), .ZN(new_n772));
  INV_X1    g0572(.A(G150), .ZN(new_n773));
  INV_X1    g0573(.A(new_n720), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT34), .Z(new_n776));
  INV_X1    g0576(.A(G132), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n708), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n722), .A2(new_n211), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n778), .B(new_n779), .C1(G58), .C2(new_n716), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n780), .B(new_n691), .C1(new_n202), .C2(new_n730), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n769), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n688), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n688), .A2(new_n682), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n702), .B1(new_n217), .B2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n783), .B(new_n785), .C1(new_n759), .C2(new_n683), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n762), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G384));
  INV_X1    g0588(.A(KEYINPUT98), .ZN(new_n789));
  INV_X1    g0589(.A(new_n397), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n399), .A2(new_n404), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT76), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n404), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n317), .B1(new_n795), .B2(KEYINPUT16), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n411), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n416), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n789), .B1(new_n799), .B2(new_n617), .ZN(new_n800));
  INV_X1    g0600(.A(new_n411), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n407), .B(new_n295), .C1(new_n795), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n417), .ZN(new_n803));
  INV_X1    g0603(.A(new_n617), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n803), .A2(KEYINPUT98), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n433), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n395), .B1(new_n802), .B2(new_n417), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n423), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n809), .A2(new_n800), .A3(new_n805), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT99), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT37), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n423), .A2(new_n418), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT37), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n413), .A2(new_n417), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n804), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n811), .B1(new_n810), .B2(KEYINPUT37), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n807), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT100), .ZN(new_n823));
  OAI211_X1 g0623(.A(KEYINPUT38), .B(new_n807), .C1(new_n818), .C2(new_n819), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n375), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n370), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n366), .A2(new_n620), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n368), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n377), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(new_n677), .A3(new_n759), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(KEYINPUT40), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n820), .A2(KEYINPUT100), .A3(new_n821), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n825), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT101), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n419), .A2(new_n816), .A3(new_n431), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n814), .B1(new_n813), .B2(new_n816), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n817), .A3(KEYINPUT101), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n433), .A2(new_n815), .A3(new_n804), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n821), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n846), .A2(new_n824), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT40), .B1(new_n847), .B2(new_n833), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n436), .A2(new_n677), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n753), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT102), .Z(new_n853));
  INV_X1    g0653(.A(new_n832), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n611), .A2(new_n620), .A3(new_n759), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n343), .A2(new_n619), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n825), .A3(new_n835), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n577), .A2(new_n617), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n375), .A2(new_n376), .A3(new_n620), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT39), .B1(new_n846), .B2(new_n824), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n825), .A2(new_n835), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n861), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n579), .B1(new_n663), .B2(new_n435), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n853), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n853), .A2(new_n869), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(new_n206), .C2(new_n700), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n460), .B(new_n232), .C1(new_n492), .C2(KEYINPUT35), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(KEYINPUT35), .B2(new_n492), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  OAI21_X1  g0675(.A(G77), .B1(new_n740), .B2(new_n211), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n876), .A2(new_n233), .B1(G50), .B2(new_n211), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(G1), .A3(new_n297), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT97), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT103), .ZN(G367));
  OAI221_X1 g0682(.A(new_n689), .B1(new_n227), .B2(new_n319), .C1(new_n693), .C2(new_n243), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n751), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n550), .A2(new_n570), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n885), .A2(new_n620), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n594), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n651), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n705), .A2(new_n202), .B1(new_n708), .B2(new_n772), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n327), .B(new_n890), .C1(G150), .C2(new_n712), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n765), .A2(G58), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n720), .A2(new_n734), .B1(new_n723), .B2(G77), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n715), .A2(new_n211), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(G143), .B2(new_n718), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n712), .A2(G303), .B1(new_n733), .B2(G317), .ZN(new_n897));
  INV_X1    g0697(.A(G283), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n705), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n447), .A2(new_n774), .B1(new_n771), .B2(new_n706), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n715), .A2(new_n328), .B1(new_n722), .B2(new_n350), .ZN(new_n901));
  OR4_X1    g0701(.A1(new_n691), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n730), .A2(new_n460), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT46), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n896), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT107), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT47), .Z(new_n907));
  INV_X1    g0707(.A(new_n688), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n884), .B1(new_n685), .B2(new_n889), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n701), .B(KEYINPUT106), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n595), .A2(new_n619), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n517), .B(new_n520), .C1(new_n518), .C2(new_n620), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n641), .A2(new_n639), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT45), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n641), .A2(new_n639), .ZN(new_n918));
  INV_X1    g0718(.A(new_n914), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT44), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n918), .A2(KEYINPUT44), .A3(new_n919), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n750), .A3(new_n637), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n638), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n641), .B1(new_n637), .B2(new_n640), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n749), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n680), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n644), .B(KEYINPUT41), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n911), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT105), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n641), .B2(new_n919), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n484), .A2(KEYINPUT105), .A3(new_n640), .A4(new_n914), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(KEYINPUT42), .A3(new_n934), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n517), .B1(new_n913), .B2(new_n483), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n937), .A2(new_n938), .B1(new_n620), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT43), .B1(new_n889), .B2(KEYINPUT104), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n940), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n638), .A2(new_n919), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n909), .B1(new_n931), .B2(new_n950), .ZN(G387));
  NOR2_X1   g0751(.A1(new_n679), .A2(new_n927), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n644), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n749), .B(new_n926), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n680), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(KEYINPUT108), .A3(new_n911), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n927), .B2(new_n910), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n634), .A2(new_n636), .A3(new_n686), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n643), .A2(new_n695), .B1(G107), .B2(new_n227), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n240), .A2(new_n272), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT109), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n643), .B(new_n272), .C1(new_n211), .C2(new_n217), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n286), .A2(new_n202), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT50), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(KEYINPUT110), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n693), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n960), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n689), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n751), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n715), .A2(new_n319), .ZN(new_n973));
  INV_X1    g0773(.A(new_n286), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n774), .A2(new_n974), .B1(new_n350), .B2(new_n722), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G159), .C2(new_n718), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n711), .A2(new_n202), .B1(new_n705), .B2(new_n211), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G150), .B2(new_n733), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n765), .A2(G77), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n976), .A2(new_n691), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n730), .A2(new_n447), .B1(new_n898), .B2(new_n715), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n712), .A2(G317), .B1(new_n742), .B2(G303), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n718), .A2(G322), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n706), .C2(new_n774), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT48), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n985), .B2(new_n984), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT49), .Z(new_n988));
  NAND2_X1  g0788(.A1(new_n723), .A2(G116), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n733), .A2(G326), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n692), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n980), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n972), .B1(new_n992), .B2(new_n688), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n956), .A2(new_n958), .B1(new_n959), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n955), .A2(new_n994), .ZN(G393));
  XNOR2_X1  g0795(.A(new_n922), .B(new_n638), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n644), .B1(new_n996), .B2(new_n952), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n925), .B1(new_n679), .B2(new_n927), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n911), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n689), .B1(new_n350), .B2(new_n227), .C1(new_n693), .C2(new_n247), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n702), .B1(new_n1001), .B2(KEYINPUT111), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT111), .B2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G317), .A2(new_n718), .B1(new_n712), .B2(G311), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT52), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n765), .A2(G283), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n327), .B1(new_n705), .B2(new_n447), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G322), .B2(new_n733), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n774), .A2(new_n731), .B1(new_n722), .B2(new_n219), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G116), .B2(new_n716), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(G143), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n722), .A2(new_n213), .B1(new_n708), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1013), .B(new_n692), .C1(new_n765), .C2(G68), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT113), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G150), .A2(new_n718), .B1(new_n712), .B2(G159), .ZN(new_n1016));
  XOR2_X1   g0816(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1017));
  XOR2_X1   g0817(.A(new_n1016), .B(new_n1017), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n716), .A2(G77), .B1(new_n742), .B2(new_n286), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n202), .C2(new_n774), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1011), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1003), .B1(new_n1021), .B2(new_n688), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n914), .B2(new_n685), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n999), .A2(new_n1000), .A3(new_n1023), .ZN(G390));
  AOI21_X1  g0824(.A(new_n702), .B1(new_n974), .B2(new_n784), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n730), .A2(new_n773), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT53), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n327), .B1(new_n733), .B2(G125), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G159), .A2(new_n716), .B1(new_n720), .B2(G137), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT54), .B(G143), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n712), .A2(G132), .B1(new_n742), .B2(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n718), .A2(G128), .B1(new_n723), .B2(G50), .ZN(new_n1033));
  AND4_X1   g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT115), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n718), .A2(G283), .B1(new_n742), .B2(G97), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n328), .B2(new_n774), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT116), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n327), .B1(new_n708), .B2(new_n447), .C1(new_n711), .C2(new_n460), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n779), .B(new_n1041), .C1(G77), .C2(new_n716), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n213), .C2(new_n730), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1027), .A2(KEYINPUT115), .A3(new_n1034), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1025), .B1(new_n908), .B2(new_n1045), .C1(new_n866), .C2(new_n683), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n832), .A2(new_n677), .A3(G330), .A4(new_n759), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n858), .A2(new_n863), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n824), .A2(new_n823), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n810), .A2(KEYINPUT37), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT99), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n817), .A3(new_n812), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT38), .B1(new_n1055), .B2(new_n807), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n835), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT39), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n864), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1051), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n759), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n857), .B1(new_n659), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n863), .B1(new_n1064), .B2(new_n832), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n846), .A2(new_n824), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1050), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT39), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n825), .B2(new_n835), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1071), .A2(new_n864), .B1(new_n863), .B2(new_n858), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n1049), .A3(new_n1067), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n644), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n677), .A2(G330), .A3(new_n759), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n854), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n856), .B1(new_n655), .B2(new_n759), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1078), .A2(new_n1047), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n856), .B1(new_n662), .B2(new_n759), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1078), .B2(new_n1047), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n379), .A2(G330), .A3(new_n434), .A4(new_n677), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n579), .B(new_n1085), .C1(new_n663), .C2(new_n435), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1076), .B1(new_n1074), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1046), .B1(new_n1075), .B2(new_n910), .C1(new_n1090), .C2(new_n1091), .ZN(G378));
  XOR2_X1   g0892(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n303), .A2(new_n804), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT55), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n310), .A2(new_n313), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n310), .B2(new_n313), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1099), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n682), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n765), .A2(new_n1031), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n711), .A2(new_n1108), .B1(new_n705), .B2(new_n772), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G125), .B2(new_n718), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G150), .A2(new_n716), .B1(new_n720), .B2(G132), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n723), .A2(new_n734), .ZN(new_n1114));
  AOI211_X1 g0914(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G41), .B1(new_n691), .B2(G33), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(G50), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n771), .A2(new_n460), .B1(new_n722), .B2(new_n740), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n894), .B(new_n1121), .C1(G97), .C2(new_n720), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n711), .A2(new_n219), .B1(new_n708), .B2(new_n898), .ZN(new_n1123));
  AOI211_X1 g0923(.A(G41), .B(new_n1123), .C1(new_n320), .C2(new_n742), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1122), .A2(new_n1124), .A3(new_n692), .A4(new_n979), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT58), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1120), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1126), .B2(new_n1125), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n688), .B1(new_n1118), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT118), .Z(new_n1130));
  AOI21_X1  g0930(.A(new_n702), .B1(new_n202), .B2(new_n784), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT119), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1104), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n849), .A2(G330), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1103), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1103), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n849), .A2(new_n1137), .A3(G330), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n867), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n861), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1059), .A2(new_n863), .A3(new_n1060), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1137), .B1(new_n849), .B2(G330), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n753), .B(new_n1103), .C1(new_n836), .C2(new_n848), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1134), .B1(new_n1146), .B2(new_n911), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1139), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1142), .B(KEYINPUT121), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT57), .B1(new_n1091), .B2(new_n1086), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1076), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1061), .A2(new_n1050), .A3(new_n1068), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1049), .B1(new_n1072), .B2(new_n1067), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1089), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1087), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT57), .B1(new_n1157), .B2(new_n1146), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1147), .B1(new_n1153), .B2(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1088), .A2(new_n930), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n702), .B1(new_n211), .B2(new_n784), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n712), .A2(G137), .B1(new_n742), .B2(G150), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1108), .B2(new_n708), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n777), .A2(new_n771), .B1(new_n774), .B2(new_n1030), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n715), .A2(new_n202), .B1(new_n722), .B2(new_n740), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n692), .B1(new_n765), .B2(G159), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n257), .B1(new_n329), .B2(new_n742), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n973), .B1(G77), .B2(new_n723), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n712), .A2(G283), .B1(new_n733), .B2(G303), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G116), .A2(new_n720), .B1(new_n718), .B2(G294), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n765), .A2(G97), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1167), .A2(new_n1168), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1162), .B1(new_n908), .B2(new_n1175), .C1(new_n832), .C2(new_n683), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1083), .B2(new_n910), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1161), .A2(new_n1178), .ZN(G381));
  NAND3_X1  g0979(.A1(new_n955), .A2(new_n755), .A3(new_n994), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1180), .A2(G381), .A3(G384), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1000), .A2(new_n1023), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n998), .B2(new_n997), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n909), .C1(new_n931), .C2(new_n950), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(G375), .A2(G378), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1187), .A2(new_n1188), .ZN(G407));
  NAND2_X1  g0989(.A1(new_n618), .A2(G213), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT123), .Z(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G407), .B(G213), .C1(new_n1188), .C2(new_n1192), .ZN(G409));
  OAI211_X1 g0993(.A(G378), .B(new_n1147), .C1(new_n1153), .C2(new_n1158), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1157), .A2(new_n930), .A3(new_n1146), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1149), .A2(new_n911), .A3(new_n1150), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1195), .A2(new_n1196), .A3(new_n1133), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1046), .B1(new_n1075), .B2(new_n910), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1194), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1083), .A2(new_n1086), .A3(KEYINPUT60), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1203), .A2(new_n1076), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1160), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G384), .B1(new_n1207), .B2(new_n1178), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1177), .B(new_n787), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1202), .A2(new_n1190), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT63), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(G387), .A2(G390), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1184), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT127), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1180), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1184), .A2(new_n1214), .A3(KEYINPUT127), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1180), .A3(new_n1218), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT61), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1202), .A2(new_n1190), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  XOR2_X1   g1027(.A(KEYINPUT124), .B(G2897), .Z(new_n1228));
  NAND3_X1  g1028(.A1(new_n618), .A2(new_n1228), .A3(G213), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1210), .B2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n618), .A2(new_n1228), .A3(G213), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1208), .A2(new_n1209), .A3(KEYINPUT125), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1191), .A2(G2897), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1230), .A2(new_n1232), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1226), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1191), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(KEYINPUT63), .A3(new_n1210), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1213), .A2(new_n1225), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1237), .B2(new_n1234), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT62), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1211), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(KEYINPUT62), .A3(new_n1210), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1241), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1224), .A2(new_n1221), .A3(new_n1220), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1239), .B1(new_n1245), .B2(new_n1247), .ZN(G405));
  NAND2_X1  g1048(.A1(G375), .A2(new_n1200), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1194), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1210), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1249), .B(new_n1194), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1246), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1246), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G402));
endmodule


