//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n206), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n211), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n221), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n214), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n247), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n225), .B1(new_n210), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n226), .A2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(G50), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n226), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n226), .B1(new_n201), .B2(new_n202), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n254), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n260), .B(new_n268), .C1(G50), .C2(new_n252), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT72), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT10), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G1698), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G1698), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G222), .B1(G77), .B2(new_n283), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n274), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n274), .A2(G274), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n274), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n286), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G200), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n271), .A2(new_n272), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n270), .A3(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n269), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n256), .A2(new_n203), .A3(new_n258), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n264), .B1(G20), .B2(G77), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n262), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n255), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n252), .A2(G77), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n297), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n289), .B1(new_n324), .B2(G244), .ZN(new_n325));
  XOR2_X1   g0125(.A(new_n325), .B(KEYINPUT70), .Z(new_n326));
  INV_X1    g0126(.A(new_n274), .ZN(new_n327));
  INV_X1    g0127(.A(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n275), .A2(new_n328), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n329), .A2(KEYINPUT71), .A3(new_n214), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT71), .B1(new_n329), .B2(new_n214), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n207), .C2(new_n275), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n277), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n327), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n323), .B1(new_n336), .B2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n336), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n310), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n326), .A2(new_n335), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n322), .B1(new_n341), .B2(new_n308), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(G58), .B2(G68), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n275), .A2(new_n350), .A3(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n283), .B2(new_n226), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n349), .B(KEYINPUT16), .C1(new_n353), .C2(new_n354), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(new_n254), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n256), .A2(new_n261), .A3(new_n258), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n250), .A2(new_n251), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n261), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n364), .B1(new_n329), .B2(new_n278), .C1(new_n298), .C2(new_n276), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n327), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n289), .B1(new_n324), .B2(G232), .ZN(new_n367));
  AOI21_X1  g0167(.A(G169), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n370), .B2(new_n310), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT18), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n363), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n370), .A2(G190), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n369), .A2(G200), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n359), .A3(new_n362), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n344), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT73), .B1(new_n253), .B2(new_n206), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT73), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(G33), .A3(G97), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G226), .A2(G1698), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n214), .B2(G1698), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n275), .B2(new_n387), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n290), .B1(new_n297), .B2(new_n333), .C1(new_n388), .C2(new_n274), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT13), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT14), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(G169), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n310), .B2(new_n390), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n390), .B2(G169), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n252), .A2(G68), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT12), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n354), .A2(G20), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(new_n262), .B2(new_n203), .C1(new_n265), .C2(new_n202), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n254), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT11), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n257), .A2(G68), .A3(new_n259), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n393), .A2(new_n394), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n390), .A2(G200), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n402), .A2(new_n396), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n404), .B(new_n405), .C1(new_n406), .C2(new_n390), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n313), .A2(new_n381), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n292), .A2(G1), .ZN(new_n410));
  AND2_X1   g0210(.A1(KEYINPUT5), .A2(G41), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT5), .A2(G41), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n287), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT5), .B(G41), .ZN(new_n415));
  INV_X1    g0215(.A(new_n225), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n415), .A2(new_n410), .B1(new_n416), .B2(new_n273), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT84), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(G264), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(G264), .A3(new_n274), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT84), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(G1698), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(new_n328), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G294), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT83), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT83), .A4(new_n425), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n406), .B(new_n422), .C1(new_n430), .C2(new_n274), .ZN(new_n431));
  INV_X1    g0231(.A(new_n414), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n418), .B1(new_n417), .B2(G264), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n420), .A2(KEYINPUT84), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n274), .B1(new_n428), .B2(new_n429), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n338), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n361), .A2(new_n207), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n253), .A2(G1), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n256), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G107), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n280), .A2(new_n282), .A3(new_n226), .A4(G87), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n275), .A2(new_n450), .A3(new_n226), .A4(G87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n453), .A2(G20), .B1(new_n454), .B2(new_n207), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n207), .A3(G20), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n207), .A3(KEYINPUT80), .A4(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT24), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n447), .B1(new_n465), .B2(new_n254), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n452), .A2(new_n463), .A3(new_n460), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n463), .B1(new_n452), .B2(new_n460), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n447), .B(new_n254), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n438), .B(new_n446), .C1(new_n466), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n254), .B1(new_n467), .B2(new_n468), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n445), .B1(new_n475), .B2(new_n469), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT85), .A3(new_n438), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n476), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n435), .A2(new_n436), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G169), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n310), .B2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT86), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT86), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n414), .B1(G270), .B2(new_n417), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n275), .A2(G264), .A3(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n283), .A2(G303), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n490), .B(new_n491), .C1(new_n329), .C2(new_n215), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT77), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n492), .A2(new_n493), .A3(new_n327), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n492), .B2(new_n327), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT78), .B(new_n489), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n252), .A2(G116), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n443), .B2(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(new_n226), .C1(G33), .C2(new_n206), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n254), .C1(new_n226), .C2(G116), .ZN(new_n504));
  XOR2_X1   g0304(.A(new_n504), .B(KEYINPUT20), .Z(new_n505));
  AOI21_X1  g0305(.A(new_n308), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n498), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT21), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n498), .A2(new_n509), .A3(new_n499), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(new_n505), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G179), .B(new_n489), .C1(new_n494), .C2(new_n495), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT79), .ZN(new_n515));
  OR3_X1    g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n498), .A2(new_n499), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n512), .B1(new_n520), .B2(G190), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n338), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(G107), .B1(new_n351), .B2(new_n352), .ZN(new_n523));
  XNOR2_X1  g0323(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n206), .A2(G107), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n208), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(G20), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n264), .A2(G77), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n254), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n361), .A2(new_n206), .ZN(new_n533));
  INV_X1    g0333(.A(new_n442), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n252), .A2(new_n255), .A3(G97), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n413), .A2(G257), .A3(new_n274), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(new_n328), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n328), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n502), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n539), .B1(new_n545), .B2(new_n327), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n546), .A2(G179), .A3(new_n432), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n308), .B1(new_n546), .B2(new_n432), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n538), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n536), .B1(new_n531), .B2(new_n254), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(G190), .A3(new_n432), .ZN(new_n551));
  AOI211_X1 g0351(.A(new_n414), .B(new_n539), .C1(new_n545), .C2(new_n327), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n338), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n317), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n443), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n252), .A2(new_n555), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n275), .A2(new_n226), .A3(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n262), .B2(new_n206), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G87), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n206), .A3(new_n207), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n560), .B1(new_n382), .B2(new_n384), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G20), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n556), .B(new_n558), .C1(new_n567), .C2(new_n255), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n274), .B(G250), .C1(G1), .C2(new_n292), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n274), .A2(G274), .A3(new_n410), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n329), .A2(new_n333), .B1(new_n253), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n275), .A2(KEYINPUT76), .A3(G244), .A4(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n310), .B(new_n572), .C1(new_n579), .C2(new_n274), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n284), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n274), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n571), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n568), .B(new_n580), .C1(new_n584), .C2(G169), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n583), .B2(new_n571), .ZN(new_n586));
  OAI211_X1 g0386(.A(G190), .B(new_n572), .C1(new_n579), .C2(new_n274), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n255), .B1(new_n562), .B2(new_n566), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n256), .A2(new_n563), .A3(new_n442), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(new_n557), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n554), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n519), .A2(new_n522), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n409), .A2(new_n488), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(G372));
  INV_X1    g0395(.A(new_n312), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n340), .A2(new_n342), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n407), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n403), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(KEYINPUT92), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT17), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n379), .B(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n599), .B2(KEYINPUT92), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n376), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n596), .B1(new_n605), .B2(new_n307), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n571), .A2(KEYINPUT87), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n569), .A2(new_n608), .A3(new_n570), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n308), .B1(new_n583), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n568), .A3(new_n580), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n583), .B2(new_n610), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n587), .A3(new_n590), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n549), .A2(new_n553), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n475), .A2(new_n469), .ZN(new_n617));
  AND4_X1   g0417(.A1(KEYINPUT85), .A2(new_n617), .A3(new_n446), .A4(new_n438), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT85), .B1(new_n476), .B2(new_n438), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n478), .A2(KEYINPUT88), .A3(new_n616), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n511), .A2(new_n483), .A3(new_n518), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT89), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT88), .B1(new_n478), .B2(new_n616), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n621), .B(new_n615), .C1(new_n473), .C2(new_n477), .ZN(new_n628));
  OAI211_X1 g0428(.A(KEYINPUT89), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  INV_X1    g0430(.A(new_n612), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n546), .A2(G179), .A3(new_n432), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n552), .B2(new_n308), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n585), .A2(new_n591), .A3(new_n633), .A4(new_n538), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n634), .B2(KEYINPUT26), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n612), .A2(new_n614), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT90), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n550), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n632), .B(KEYINPUT90), .C1(new_n308), .C2(new_n552), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n636), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n630), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n635), .A2(new_n641), .A3(new_n630), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n629), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n409), .B1(new_n626), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n606), .A2(new_n647), .ZN(G369));
  INV_X1    g0448(.A(new_n487), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n486), .B1(new_n478), .B2(new_n483), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n247), .A2(new_n226), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n649), .A2(new_n650), .B1(new_n476), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n479), .A2(new_n482), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n519), .B(new_n522), .C1(new_n513), .C2(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n511), .A2(new_n518), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n513), .A2(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n661), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n657), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n485), .B2(new_n487), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n483), .A2(new_n656), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n222), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n564), .A2(G116), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n674), .A2(new_n247), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n229), .B2(new_n674), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  NAND3_X1  g0478(.A1(new_n625), .A2(new_n478), .A3(new_n616), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n612), .B1(new_n634), .B2(KEYINPUT26), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n636), .A2(new_n640), .A3(new_n638), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(KEYINPUT26), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n656), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n657), .B1(new_n646), .B2(new_n626), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n488), .A2(new_n593), .A3(new_n657), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n480), .A2(new_n584), .A3(new_n546), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n690), .A2(new_n691), .A3(new_n514), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n690), .B2(new_n514), .ZN(new_n693));
  INV_X1    g0493(.A(new_n480), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n583), .A2(new_n610), .ZN(new_n695));
  INV_X1    g0495(.A(new_n552), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n694), .A2(new_n695), .A3(new_n310), .A4(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n692), .B(new_n693), .C1(new_n520), .C2(new_n697), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT31), .B1(new_n698), .B2(new_n656), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT93), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n656), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n656), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n689), .A2(new_n701), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n688), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n678), .B1(new_n711), .B2(G1), .ZN(G364));
  AND2_X1   g0512(.A1(new_n226), .A2(G13), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n247), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n674), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n666), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n662), .A2(new_n661), .A3(new_n665), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n662), .A2(new_n665), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n225), .B1(G20), .B2(new_n308), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n722), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n222), .A2(new_n275), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT94), .Z(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n573), .B2(new_n673), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n242), .A2(G45), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n673), .A2(new_n275), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n734), .C1(G45), .C2(new_n228), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n729), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n727), .ZN(new_n737));
  NAND2_X1  g0537(.A1(G20), .A2(G179), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G190), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n738), .A2(new_n406), .A3(G200), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n742), .A2(G77), .B1(G58), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n738), .A2(new_n338), .A3(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n354), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n226), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n740), .ZN(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n753), .A2(KEYINPUT32), .A3(G159), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n747), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n226), .A2(new_n338), .A3(G179), .A4(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n406), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n226), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n757), .A2(new_n207), .B1(new_n759), .B2(new_n206), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n739), .A2(G190), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(G50), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n275), .B1(new_n764), .B2(new_n563), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n755), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  INV_X1    g0568(.A(G294), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n757), .A2(new_n768), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n745), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n750), .B(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  INV_X1    g0574(.A(new_n743), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n283), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G311), .B2(new_n742), .ZN(new_n778));
  INV_X1    g0578(.A(new_n764), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G303), .A2(new_n779), .B1(new_n762), .B2(G326), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n772), .A2(new_n774), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n737), .B1(new_n767), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n716), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n736), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n723), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n719), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  OAI211_X1 g0587(.A(new_n344), .B(new_n657), .C1(new_n646), .C2(new_n626), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n635), .A2(new_n641), .A3(new_n630), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n642), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n511), .A2(new_n483), .A3(new_n518), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n622), .B2(new_n623), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(KEYINPUT89), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT89), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n656), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n343), .A2(new_n656), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n323), .A2(new_n656), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n339), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n800), .B2(new_n343), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n788), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(new_n709), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n716), .B1(new_n802), .B2(new_n709), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n283), .B1(new_n779), .B2(G50), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n213), .B2(new_n759), .C1(new_n354), .C2(new_n757), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n742), .A2(G159), .B1(G143), .B2(new_n743), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n263), .B2(new_n746), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G137), .B2(new_n762), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n807), .B(new_n811), .C1(G132), .C2(new_n773), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n773), .A2(G311), .B1(G87), .B2(new_n756), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT99), .Z(new_n814));
  OAI221_X1 g0614(.A(new_n283), .B1(new_n741), .B2(new_n573), .C1(new_n775), .C2(new_n769), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n759), .A2(new_n206), .B1(new_n746), .B2(new_n768), .ZN(new_n816));
  INV_X1    g0616(.A(G303), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n764), .A2(new_n207), .B1(new_n761), .B2(new_n817), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n727), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n727), .A2(new_n720), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n716), .B1(new_n822), .B2(G77), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT98), .Z(new_n824));
  OAI211_X1 g0624(.A(new_n820), .B(new_n824), .C1(new_n801), .C2(new_n721), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n805), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  NAND2_X1  g0628(.A1(new_n526), .A2(new_n528), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT35), .ZN(new_n830));
  OAI211_X1 g0630(.A(G116), .B(new_n227), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n347), .A2(G77), .A3(new_n229), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n202), .A2(G68), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n247), .B(G13), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n798), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n788), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n654), .B1(new_n359), .B2(new_n362), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT101), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n373), .A2(new_n375), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n842), .B(new_n844), .C1(new_n602), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n844), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n372), .A2(new_n379), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n840), .A3(KEYINPUT37), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n846), .B(KEYINPUT38), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n405), .B(new_n657), .C1(new_n403), .C2(new_n407), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n405), .A2(new_n657), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n408), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n839), .A2(new_n857), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n845), .A2(new_n654), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n847), .B1(new_n850), .B2(new_n841), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n852), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n841), .B1(new_n376), .B2(new_n380), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n854), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n856), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g0671(.A1(new_n403), .A2(KEYINPUT102), .A3(new_n656), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT102), .B1(new_n403), .B2(new_n656), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n863), .A2(new_n864), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n845), .B1(new_n600), .B2(new_n603), .ZN(new_n878));
  INV_X1    g0678(.A(new_n307), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n312), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n688), .B2(new_n409), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n877), .B(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n699), .A2(new_n700), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n689), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n801), .B1(new_n858), .B2(new_n860), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n869), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT40), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT40), .B1(new_n855), .B2(new_n856), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n689), .B2(new_n883), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n409), .A2(new_n884), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n661), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n882), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n247), .B2(new_n713), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n882), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n837), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT103), .ZN(G367));
  INV_X1    g0700(.A(new_n734), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n728), .B1(new_n222), .B2(new_n317), .C1(new_n901), .C2(new_n237), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n716), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n746), .A2(new_n751), .B1(new_n764), .B2(new_n213), .ZN(new_n904));
  INV_X1    g0704(.A(new_n759), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(G68), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n283), .B1(new_n753), .B2(G137), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n742), .A2(G50), .B1(G150), .B2(new_n743), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n762), .A2(G143), .B1(new_n756), .B2(G77), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(G317), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n283), .B1(new_n911), .B2(new_n750), .C1(new_n757), .C2(new_n206), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT106), .Z(new_n913));
  INV_X1    g0713(.A(KEYINPUT46), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n764), .A2(new_n914), .A3(new_n573), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n775), .A2(new_n817), .B1(new_n741), .B2(new_n768), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G294), .B2(new_n745), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n914), .B1(new_n764), .B2(new_n573), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n905), .A2(G107), .B1(new_n762), .B2(G311), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n910), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT47), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(new_n727), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n924), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n903), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n590), .A2(new_n657), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n636), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n929), .A2(new_n612), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n722), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT104), .ZN(new_n936));
  INV_X1    g0736(.A(new_n711), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n554), .B1(new_n550), .B2(new_n657), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n638), .A2(new_n640), .A3(new_n656), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n938), .B1(new_n671), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n668), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n649), .B2(new_n650), .ZN(new_n944));
  INV_X1    g0744(.A(new_n670), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n941), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n949), .A2(new_n953), .A3(new_n667), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n667), .B1(new_n949), .B2(new_n953), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n944), .B1(new_n660), .B2(new_n943), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n666), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n937), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n674), .B(KEYINPUT41), .Z(new_n960));
  OAI21_X1  g0760(.A(new_n714), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n549), .A2(new_n656), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n669), .A2(new_n941), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n963), .B2(KEYINPUT42), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n947), .B1(KEYINPUT42), .B2(new_n945), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n946), .A2(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n964), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n667), .A2(new_n947), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n970), .A3(new_n933), .A4(new_n966), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n936), .B1(new_n961), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n671), .B2(new_n941), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT44), .B1(new_n946), .B2(new_n947), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n938), .B(new_n941), .C1(new_n944), .C2(new_n945), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n667), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n949), .A2(new_n953), .A3(new_n667), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n982), .A2(new_n711), .A3(new_n958), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n960), .B1(new_n984), .B2(new_n711), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n974), .B(new_n936), .C1(new_n985), .C2(new_n715), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n935), .B1(new_n975), .B2(new_n987), .ZN(G387));
  NAND2_X1  g0788(.A1(new_n731), .A2(new_n675), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(G107), .B2(new_n222), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n234), .A2(new_n292), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n261), .A2(G50), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  AOI211_X1 g0793(.A(G45), .B(new_n675), .C1(G68), .C2(G77), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n901), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n990), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n716), .B1(new_n996), .B2(new_n729), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n750), .A2(new_n263), .B1(new_n741), .B2(new_n354), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n283), .B(new_n998), .C1(G50), .C2(new_n743), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n779), .A2(G77), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n905), .A2(new_n555), .B1(new_n315), .B2(new_n745), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n762), .A2(G159), .B1(new_n756), .B2(G97), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n759), .A2(new_n768), .B1(new_n764), .B2(new_n769), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n742), .A2(G303), .B1(G317), .B2(new_n743), .ZN(new_n1005));
  INV_X1    g0805(.A(G311), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n746), .C1(new_n776), .C2(new_n761), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n275), .B1(new_n753), .B2(G326), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n573), .B2(new_n757), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT107), .Z(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1003), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n997), .B1(new_n727), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n722), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n660), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT108), .Z(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n715), .B2(new_n958), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n958), .A2(new_n711), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n674), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n958), .A2(new_n711), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G393));
  AOI22_X1  g0826(.A1(new_n762), .A2(G317), .B1(G311), .B2(new_n743), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT52), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n283), .B1(new_n741), .B2(new_n769), .C1(new_n776), .C2(new_n750), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n757), .A2(new_n207), .B1(new_n817), .B2(new_n746), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n759), .A2(new_n573), .B1(new_n764), .B2(new_n768), .ZN(new_n1031));
  OR4_X1    g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n759), .A2(new_n203), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n746), .A2(new_n202), .B1(new_n764), .B2(new_n354), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G87), .C2(new_n756), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n775), .A2(new_n751), .B1(new_n761), .B2(new_n263), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n753), .A2(G143), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n283), .B1(new_n742), .B2(new_n315), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n737), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n734), .A2(new_n245), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n729), .B1(G97), .B2(new_n673), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n783), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n941), .B2(new_n1019), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n982), .A2(new_n983), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n714), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n984), .A2(new_n674), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1023), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G390));
  NAND2_X1  g0851(.A1(new_n871), .A2(new_n875), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n861), .B1(new_n788), .B2(new_n838), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n874), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n661), .B1(new_n689), .B2(new_n883), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(KEYINPUT110), .A3(new_n886), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n710), .A2(new_n1056), .A3(new_n801), .A4(new_n862), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n800), .A2(new_n343), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n798), .B1(new_n683), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n862), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n874), .A2(KEYINPUT109), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n874), .A2(KEYINPUT109), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1061), .A2(new_n869), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1054), .A2(new_n1057), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1055), .A2(new_n886), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT110), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1054), .B2(new_n1064), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n409), .B(new_n684), .C1(new_n797), .C2(KEYINPUT29), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1055), .A2(new_n409), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n606), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT111), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n708), .A2(G330), .A3(new_n801), .A4(new_n862), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1058), .A2(new_n838), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n661), .B(new_n1078), .C1(new_n689), .C2(new_n883), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1077), .B(new_n1059), .C1(new_n862), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n839), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n488), .A2(new_n593), .A3(new_n657), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n701), .A2(new_n707), .ZN(new_n1083));
  OAI211_X1 g0883(.A(G330), .B(new_n801), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1084), .A2(new_n861), .B1(new_n886), .B2(new_n1055), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1080), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1072), .A2(new_n606), .A3(KEYINPUT111), .A4(new_n1073), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1076), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(KEYINPUT112), .B1(new_n1071), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n674), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1071), .B2(new_n1088), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1076), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT112), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n1065), .C2(new_n1070), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n275), .B1(new_n757), .B2(new_n202), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1096), .A2(new_n1097), .B1(new_n773), .B2(G125), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT115), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n779), .A2(G150), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n905), .A2(G159), .B1(G137), .B2(new_n745), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n762), .A2(G128), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n742), .A2(new_n1106), .B1(G132), .B2(new_n743), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1100), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n761), .A2(new_n768), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1033), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n207), .B2(new_n746), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n773), .A2(G294), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n283), .B1(new_n741), .B2(new_n206), .C1(new_n775), .C2(new_n573), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n757), .A2(new_n354), .B1(new_n563), .B2(new_n764), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n727), .B1(new_n1109), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n716), .C1(new_n315), .C2(new_n822), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1052), .B2(new_n720), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1054), .A2(new_n1057), .A3(new_n1064), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1054), .A2(new_n1064), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n715), .B(new_n1120), .C1(new_n1121), .C2(new_n1069), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT113), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1070), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n715), .A4(new_n1120), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1119), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1095), .A2(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1076), .A2(new_n1087), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1071), .B2(new_n1088), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n654), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n269), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n313), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n313), .A2(new_n1136), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1137), .A3(new_n1132), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n892), .A2(G330), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n887), .A2(KEYINPUT40), .B1(new_n889), .B2(new_n890), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n661), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n877), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n877), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1129), .B1(new_n1131), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n877), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1148), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1092), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(KEYINPUT57), .C1(new_n1157), .C2(new_n1130), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n674), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n715), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n283), .A2(new_n291), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n779), .B2(G77), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n213), .B2(new_n757), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G283), .B2(new_n773), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT116), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n775), .A2(new_n207), .B1(new_n317), .B2(new_n741), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G68), .B2(new_n905), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n762), .A2(G116), .B1(G97), .B2(new_n745), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1161), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1171));
  INV_X1    g0971(.A(G132), .ZN(new_n1172));
  INV_X1    g0972(.A(G125), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n746), .A2(new_n1172), .B1(new_n761), .B2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n742), .A2(G137), .B1(G128), .B2(new_n743), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n764), .B2(new_n1105), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G150), .C2(new_n905), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT117), .Z(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(KEYINPUT59), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n751), .B2(new_n757), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT118), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1170), .B(new_n1171), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT119), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n727), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT120), .Z(new_n1189));
  AOI21_X1  g0989(.A(new_n783), .B1(new_n202), .B2(new_n821), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n721), .C2(new_n1143), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1160), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1159), .A2(new_n1193), .ZN(G375));
  NAND2_X1  g0994(.A1(new_n1084), .A2(new_n861), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1066), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1055), .A2(new_n801), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1060), .B1(new_n1197), .B2(new_n861), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1196), .A2(new_n839), .B1(new_n1198), .B2(new_n1077), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT111), .B1(new_n881), .B2(new_n1073), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1087), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1086), .B1(new_n1076), .B2(new_n1087), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT121), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n960), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .A4(new_n1092), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n861), .A2(new_n720), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n764), .A2(new_n206), .B1(new_n761), .B2(new_n769), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G116), .B2(new_n745), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n773), .A2(G303), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n283), .B1(new_n741), .B2(new_n207), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n743), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n905), .A2(new_n555), .B1(G77), .B2(new_n756), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n764), .A2(new_n751), .B1(new_n761), .B2(new_n1172), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G50), .B2(new_n905), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n773), .A2(G128), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n275), .B1(new_n741), .B2(new_n263), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G137), .B2(new_n743), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n745), .A2(new_n1106), .B1(new_n756), .B2(G58), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n737), .B1(new_n1216), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n783), .B(new_n1224), .C1(new_n354), .C2(new_n821), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1086), .A2(new_n715), .B1(new_n1209), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1208), .A2(new_n1226), .ZN(G381));
  NAND2_X1  g1027(.A1(new_n1050), .A2(new_n827), .ZN(new_n1228));
  OR4_X1    g1028(.A1(G396), .A2(G387), .A3(G393), .A4(new_n1228), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G375), .A3(G381), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT122), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1095), .A2(new_n1127), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n1095), .B2(new_n1127), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n1234), .ZN(G407));
  NAND2_X1  g1035(.A1(new_n655), .A2(G213), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT123), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1193), .A3(new_n1159), .A4(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  INV_X1    g1039(.A(new_n1237), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1131), .A2(new_n1151), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1192), .B1(new_n1241), .B2(new_n1207), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1232), .A2(new_n1233), .A3(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1159), .A2(G378), .A3(new_n1193), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1240), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1204), .A2(new_n1206), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1090), .B1(new_n1205), .B2(KEYINPUT60), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1226), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n827), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G384), .B(new_n1226), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT62), .B1(new_n1245), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1237), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT124), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1262), .B2(new_n1226), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1254), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1253), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1245), .A3(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1095), .A2(new_n1127), .A3(new_n1231), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1156), .B1(new_n1157), .B2(new_n1130), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1193), .B1(new_n1272), .B2(new_n960), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1159), .A2(G378), .A3(new_n1193), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1237), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1269), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1256), .A2(new_n1267), .A3(new_n1268), .A4(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n786), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n974), .B1(new_n985), .B2(new_n715), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT104), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n986), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G390), .B1(new_n1284), .B2(new_n935), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n935), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1286), .B(new_n1050), .C1(new_n1283), .C2(new_n986), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G387), .A2(new_n1050), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1284), .A2(G390), .A3(new_n935), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1280), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1279), .A2(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1254), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1292), .B1(new_n1294), .B2(new_n1276), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1245), .B2(new_n1255), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1295), .A2(new_n1297), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1298), .A2(KEYINPUT125), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1254), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1245), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT63), .B1(new_n1269), .B2(new_n1276), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1257), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(new_n1276), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1266), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1300), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1293), .B1(new_n1299), .B2(new_n1309), .ZN(G405));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1234), .A2(new_n1311), .A3(G375), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1275), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1234), .B2(G375), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(KEYINPUT127), .A3(new_n1269), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1255), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1317), .B(new_n1319), .C1(new_n1314), .C2(new_n1313), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1316), .A2(new_n1301), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1301), .B1(new_n1316), .B2(new_n1320), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


