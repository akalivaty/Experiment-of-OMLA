//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT24), .B(G110), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G119), .B(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G110), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT78), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n193), .B2(G119), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n195), .A2(new_n196), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G125), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT79), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n203), .B1(new_n207), .B2(new_n199), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n202), .B1(new_n208), .B2(new_n201), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(G146), .ZN(new_n212));
  OAI221_X1 g026(.A(new_n191), .B1(new_n192), .B2(new_n198), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n198), .A2(new_n192), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n190), .B2(new_n189), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT64), .A2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n215), .B(new_n210), .C1(new_n218), .C2(new_n207), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n221), .B(new_n223), .Z(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n213), .A2(new_n219), .A3(new_n224), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G234), .B2(new_n227), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n231), .A2(KEYINPUT80), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT80), .B1(new_n231), .B2(new_n233), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n228), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n237), .A2(G902), .A3(new_n233), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n187), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NOR4_X1   g054(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT81), .A4(new_n238), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT64), .A2(G146), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT64), .A2(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(new_n251), .B2(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n252), .A2(new_n193), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n216), .A2(G143), .A3(new_n217), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(G146), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n248), .A3(G128), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G134), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(G134), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT65), .A2(G134), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT65), .A2(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n262), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n256), .A2(new_n259), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT11), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(G134), .B2(new_n261), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT65), .A2(G134), .ZN(new_n279));
  AOI21_X1  g093(.A(G137), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n275), .B1(new_n280), .B2(new_n274), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n265), .B1(new_n263), .B2(new_n261), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT66), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n274), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n284));
  INV_X1    g098(.A(new_n275), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n267), .A2(new_n268), .ZN(new_n287));
  AOI21_X1  g101(.A(G131), .B1(new_n287), .B2(G137), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n247), .B1(new_n273), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n263), .A2(new_n261), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n281), .B2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n289), .B1(new_n286), .B2(new_n288), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n255), .B1(new_n218), .B2(new_n254), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n257), .A2(new_n258), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  OAI22_X1  g115(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n292), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n222), .A3(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT27), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G101), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n193), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n259), .B1(new_n313), .B2(new_n298), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n266), .A2(new_n272), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n291), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(new_n247), .B1(new_n292), .B2(new_n304), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n307), .B(new_n312), .C1(new_n318), .C2(new_n306), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n227), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n322), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n304), .A2(new_n327), .A3(new_n316), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n304), .B2(new_n316), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n247), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n305), .ZN(new_n331));
  INV_X1    g145(.A(new_n312), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n333), .A3(new_n320), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G472), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g151(.A(new_n247), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n295), .A2(new_n296), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n271), .A2(KEYINPUT67), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n260), .B(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n314), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n338), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n302), .B1(new_n291), .B2(new_n294), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n312), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n305), .A2(KEYINPUT69), .A3(new_n312), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n339), .A2(new_n342), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT30), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n304), .A2(new_n316), .A3(new_n327), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n347), .A2(new_n348), .B1(new_n352), .B2(new_n247), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n307), .B1(new_n318), .B2(new_n306), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n332), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT70), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n347), .A2(new_n348), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n357), .B(new_n354), .C1(new_n358), .C2(new_n330), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT69), .B1(new_n305), .B2(new_n312), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n346), .B(new_n332), .C1(new_n292), .C2(new_n304), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n330), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT70), .B1(new_n362), .B2(KEYINPUT31), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n356), .C1(new_n359), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(KEYINPUT32), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n335), .A2(new_n371), .A3(G472), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n337), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT72), .B1(new_n368), .B2(new_n369), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n376));
  INV_X1    g190(.A(new_n369), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n376), .B(new_n377), .C1(new_n365), .C2(new_n367), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT73), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n367), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n357), .B1(new_n353), .B2(new_n354), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n362), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n366), .B1(new_n385), .B2(new_n356), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n369), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n376), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n368), .A2(KEYINPUT72), .A3(new_n369), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n388), .A2(KEYINPUT73), .A3(new_n380), .A4(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n374), .B1(new_n381), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n380), .A3(new_n389), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n390), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n374), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n243), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n302), .A2(G125), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(G125), .B2(new_n314), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n222), .A2(G224), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g219(.A(G104), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G107), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G104), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G101), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n410), .A2(KEYINPUT83), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT83), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n406), .C2(G107), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n409), .B1(new_n416), .B2(new_n407), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n411), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n244), .A2(KEYINPUT5), .ZN(new_n422));
  INV_X1    g236(.A(G116), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n423), .A2(KEYINPUT5), .A3(G119), .ZN(new_n424));
  INV_X1    g238(.A(G113), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n246), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n422), .A2(new_n426), .B1(new_n427), .B2(new_n244), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n414), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n419), .A2(new_n420), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G101), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n434), .A2(KEYINPUT4), .ZN(new_n435));
  INV_X1    g249(.A(new_n421), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(KEYINPUT4), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n435), .B(new_n247), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n430), .A3(new_n431), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(KEYINPUT85), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n441), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n441), .A2(new_n442), .B1(KEYINPUT86), .B2(KEYINPUT6), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n405), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n402), .A2(new_n449), .B1(KEYINPUT7), .B2(new_n404), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n403), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n439), .B(KEYINPUT8), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n414), .A2(new_n421), .ZN(new_n454));
  INV_X1    g268(.A(new_n244), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n422), .A2(KEYINPUT87), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n422), .A2(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n426), .ZN(new_n458));
  OAI221_X1 g272(.A(new_n454), .B1(new_n246), .B2(new_n455), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT88), .B1(new_n454), .B2(new_n428), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n454), .A2(KEYINPUT88), .A3(new_n428), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n453), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n452), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n446), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n446), .B2(new_n464), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n401), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n227), .ZN(new_n475));
  INV_X1    g289(.A(new_n259), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT1), .B1(new_n254), .B2(G146), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n257), .A2(new_n258), .B1(G128), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n454), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT10), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n297), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n435), .B(new_n303), .C1(new_n436), .C2(new_n437), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n454), .A2(KEYINPUT10), .A3(new_n314), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n479), .B1(new_n314), .B2(new_n454), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n486), .A2(KEYINPUT12), .A3(new_n297), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT12), .B1(new_n486), .B2(new_n297), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G140), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n222), .A2(G227), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n297), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n489), .A2(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n475), .B1(new_n497), .B2(G469), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n494), .B1(new_n487), .B2(new_n488), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n485), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n492), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n474), .A3(new_n227), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n473), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT90), .B(new_n401), .C1(new_n466), .C2(new_n467), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n470), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n406), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n308), .A2(new_n222), .A3(G214), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n254), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G131), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n207), .B(KEYINPUT91), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT19), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n207), .A2(KEYINPUT19), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT92), .B1(new_n518), .B2(new_n218), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n520), .A3(new_n251), .A4(new_n517), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT18), .A2(G131), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n512), .B(new_n523), .Z(new_n524));
  NOR2_X1   g338(.A1(new_n218), .A2(new_n207), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n515), .B2(G146), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n510), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n527), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n512), .A2(KEYINPUT17), .A3(G131), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT93), .ZN(new_n531));
  INV_X1    g345(.A(new_n212), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n532), .B(new_n210), .C1(new_n513), .C2(KEYINPUT17), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n529), .B(new_n509), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT20), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(KEYINPUT94), .A3(new_n534), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n536), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n541), .B1(new_n545), .B2(KEYINPUT20), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n529), .B1(new_n533), .B2(new_n531), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n534), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n227), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(G475), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n546), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(G234), .A2(G237), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G952), .A3(new_n222), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(G902), .A3(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G107), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT97), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n254), .A2(G128), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n193), .A2(G143), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n287), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(KEYINPUT13), .ZN(new_n570));
  OAI21_X1  g384(.A(G134), .B1(new_n566), .B2(KEYINPUT13), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n565), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G122), .ZN(new_n573));
  OR3_X1    g387(.A1(new_n573), .A2(KEYINPUT14), .A3(G116), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n423), .A2(G122), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT14), .B1(new_n573), .B2(G116), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT98), .A4(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(G107), .C1(KEYINPUT98), .C2(new_n574), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n568), .B(new_n287), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n563), .A2(new_n408), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n572), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n471), .A2(new_n232), .A3(G953), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n572), .A2(new_n582), .A3(new_n584), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G478), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT15), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n588), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n553), .A2(new_n554), .A3(new_n562), .A4(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n507), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n400), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n368), .A2(new_n227), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n242), .A2(new_n379), .A3(new_n504), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n586), .A2(new_n587), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT33), .B1(new_n584), .B2(KEYINPUT99), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n603), .B(new_n604), .Z(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n589), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(new_n589), .ZN(new_n607));
  NAND2_X1  g421(.A1(G478), .A2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n553), .B2(new_n554), .ZN(new_n611));
  INV_X1    g425(.A(new_n468), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n562), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n562), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n545), .B(KEYINPUT20), .ZN(new_n618));
  INV_X1    g432(.A(new_n552), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n619), .A3(new_n592), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n602), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(new_n236), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n220), .B(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n626), .A2(G902), .A3(new_n233), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n506), .A2(new_n628), .A3(new_n594), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n379), .A3(new_n601), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT37), .B(G110), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT100), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G12));
  INV_X1    g447(.A(new_n628), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n504), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n468), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT101), .B(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n557), .B1(new_n637), .B2(new_n559), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n620), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n398), .B1(new_n397), .B2(new_n374), .ZN(new_n640));
  AOI211_X1 g454(.A(KEYINPUT77), .B(new_n373), .C1(new_n396), .C2(new_n390), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n636), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  XOR2_X1   g457(.A(new_n638), .B(KEYINPUT39), .Z(new_n644));
  NAND2_X1  g458(.A1(new_n504), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT40), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n466), .A2(new_n467), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n554), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n593), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n401), .A2(new_n649), .A3(new_n628), .A4(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n318), .A2(new_n312), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n227), .B1(new_n353), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G472), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n370), .B(new_n657), .C1(new_n381), .C2(new_n391), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n646), .B1(new_n662), .B2(KEYINPUT103), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n654), .C1(new_n660), .C2(new_n661), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  INV_X1    g482(.A(new_n610), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n650), .B2(new_n651), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n668), .B1(new_n670), .B2(new_n638), .ZN(new_n671));
  INV_X1    g485(.A(new_n638), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n611), .A2(KEYINPUT104), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n636), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n640), .B2(new_n641), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NAND2_X1  g491(.A1(new_n502), .A2(new_n227), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n474), .A2(KEYINPUT105), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n679), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n502), .A2(new_n227), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n682), .A3(new_n472), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n243), .A2(new_n613), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n640), .B2(new_n641), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NOR2_X1   g501(.A1(new_n617), .A2(new_n620), .ZN(new_n688));
  INV_X1    g502(.A(new_n683), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n400), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT106), .B(G116), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G18));
  NOR2_X1   g508(.A1(new_n683), .A2(new_n468), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n594), .A3(new_n628), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n640), .B2(new_n641), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND2_X1  g513(.A1(new_n689), .A2(new_n562), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n700), .A2(new_n652), .A3(new_n593), .A4(new_n468), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n624), .A2(new_n238), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n356), .B1(new_n354), .B2(new_n353), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n369), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT108), .Z(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n601), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NAND3_X1  g523(.A1(new_n634), .A2(new_n601), .A3(new_n705), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT109), .ZN(new_n711));
  INV_X1    g525(.A(new_n696), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n674), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  INV_X1    g528(.A(new_n504), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n647), .A2(new_n401), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n674), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n242), .C1(new_n641), .C2(new_n640), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n674), .A2(KEYINPUT42), .A3(new_n719), .ZN(new_n724));
  INV_X1    g538(.A(new_n387), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n374), .B1(new_n725), .B2(KEYINPUT32), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n702), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT111), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n731), .B(new_n728), .C1(new_n721), .C2(new_n722), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  AND2_X1   g548(.A1(new_n719), .A2(new_n242), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n639), .B(new_n735), .C1(new_n640), .C2(new_n641), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G134), .ZN(G36));
  NAND2_X1  g551(.A1(new_n652), .A2(new_n669), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT43), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n628), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n379), .A2(new_n601), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n741), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n497), .B2(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(KEYINPUT45), .B2(new_n497), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n475), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT46), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n503), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n472), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n718), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(new_n644), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n744), .A2(new_n745), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NAND2_X1  g571(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n674), .A2(new_n243), .A3(new_n754), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n399), .A3(new_n393), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NOR2_X1   g578(.A1(new_n660), .A2(new_n661), .ZN(new_n765));
  INV_X1    g579(.A(new_n738), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n702), .A3(new_n401), .A4(new_n472), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT112), .ZN(new_n769));
  INV_X1    g583(.A(new_n680), .ZN(new_n770));
  INV_X1    g584(.A(new_n682), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT49), .Z(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n649), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n765), .A2(new_n768), .A3(new_n769), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n718), .A2(new_n683), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n765), .A2(new_n242), .A3(new_n557), .A4(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT116), .Z(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n652), .A3(new_n610), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n739), .A2(new_n556), .A3(new_n706), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n683), .A2(new_n401), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n649), .B1(new_n781), .B2(KEYINPUT115), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n782), .C1(KEYINPUT115), .C2(new_n781), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT50), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n739), .A2(new_n556), .A3(new_n683), .A4(new_n718), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n711), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n772), .A2(new_n473), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n758), .A2(new_n760), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(KEYINPUT117), .ZN(new_n789));
  INV_X1    g603(.A(new_n780), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n789), .A2(new_n718), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(KEYINPUT117), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n727), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n785), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  INV_X1    g613(.A(G952), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n800), .B(G953), .C1(new_n780), .C2(new_n712), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n778), .B2(new_n611), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n788), .A2(new_n754), .A3(new_n780), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n779), .A2(new_n804), .A3(new_n786), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n794), .B(new_n803), .C1(new_n805), .C2(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n720), .A2(new_n711), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n618), .A2(new_n593), .A3(new_n619), .A4(new_n672), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n635), .A2(new_n718), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n640), .B2(new_n641), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n736), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n470), .A2(new_n562), .A3(new_n505), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n670), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n470), .A2(new_n505), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n650), .A2(new_n651), .A3(new_n593), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n562), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n562), .A4(new_n611), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n602), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n630), .A2(new_n708), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n685), .A3(new_n698), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n400), .B1(new_n597), .B2(new_n691), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n811), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n730), .A3(new_n732), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n653), .A2(new_n612), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n634), .A2(new_n715), .A3(new_n638), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n658), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n642), .A2(new_n676), .A3(new_n713), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n642), .A2(new_n713), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n826), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT42), .B1(new_n400), .B2(new_n720), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n731), .B1(new_n839), .B2(new_n728), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n723), .A2(KEYINPUT111), .A3(new_n729), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n822), .A2(new_n685), .A3(new_n698), .ZN(new_n842));
  AOI221_X4 g656(.A(new_n243), .B1(new_n596), .B2(new_n690), .C1(new_n393), .C2(new_n399), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n841), .A3(new_n844), .A4(new_n811), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n831), .B(KEYINPUT52), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n836), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n723), .A2(new_n729), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n835), .ZN(new_n852));
  INV_X1    g666(.A(new_n825), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n833), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n806), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n775), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n854), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(G210), .A3(G902), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n444), .A2(new_n445), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(new_n405), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT55), .Z(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n800), .A2(G953), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT120), .Z(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(G51));
  AND3_X1   g686(.A1(new_n860), .A2(G902), .A3(new_n747), .ZN(new_n873));
  XNOR2_X1  g687(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n475), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n847), .A2(new_n850), .A3(new_n854), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n850), .B1(new_n847), .B2(new_n854), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n878), .B2(new_n502), .ZN(new_n879));
  INV_X1    g693(.A(new_n868), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT122), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n882));
  INV_X1    g696(.A(new_n502), .ZN(new_n883));
  INV_X1    g697(.A(new_n850), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT53), .B1(new_n826), .B2(new_n833), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n833), .A2(new_n852), .A3(new_n853), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n855), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n883), .B1(new_n888), .B2(new_n875), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n882), .B(new_n868), .C1(new_n889), .C2(new_n873), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n881), .A2(new_n890), .ZN(G54));
  AND2_X1   g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n860), .A2(G902), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n543), .ZN(new_n894));
  INV_X1    g708(.A(new_n544), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n860), .A2(G902), .A3(new_n897), .A4(new_n892), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n868), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(KEYINPUT123), .A3(new_n868), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G60));
  XNOR2_X1  g717(.A(new_n608), .B(KEYINPUT59), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n888), .A2(new_n605), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n605), .B1(new_n856), .B2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n880), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT60), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n847), .B2(new_n854), .ZN(new_n910));
  INV_X1    g724(.A(new_n626), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n237), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n868), .C1(new_n913), .C2(new_n910), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G66));
  INV_X1    g730(.A(new_n560), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n222), .B1(new_n917), .B2(G224), .ZN(new_n918));
  INV_X1    g732(.A(new_n844), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n222), .ZN(new_n920));
  INV_X1    g734(.A(G898), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n863), .B1(new_n921), .B2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n920), .B(new_n922), .ZN(G69));
  XOR2_X1   g737(.A(new_n352), .B(new_n518), .Z(new_n924));
  NAND2_X1  g738(.A1(G900), .A2(G953), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n642), .A2(new_n676), .A3(new_n713), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n795), .A2(new_n644), .A3(new_n828), .A4(new_n753), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n736), .A2(new_n756), .A3(new_n763), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n733), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT126), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n924), .B(new_n925), .C1(new_n931), .C2(G953), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n645), .A2(new_n718), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n400), .B(new_n933), .C1(new_n611), .C2(new_n816), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n763), .A3(new_n756), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n666), .A2(new_n927), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(KEYINPUT62), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n926), .B1(new_n663), .B2(new_n665), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n938), .A2(KEYINPUT124), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT125), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n937), .B(new_n944), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  AOI21_X1  g759(.A(G953), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n932), .B1(new_n946), .B2(new_n924), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n932), .B(new_n950), .C1(new_n946), .C2(new_n924), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G72));
  XOR2_X1   g766(.A(new_n331), .B(KEYINPUT127), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n844), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI211_X1 g770(.A(new_n332), .B(new_n953), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n333), .B2(new_n362), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n880), .B1(new_n848), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n931), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n961), .B2(new_n844), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n953), .A2(new_n332), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n957), .A2(new_n964), .ZN(G57));
endmodule


