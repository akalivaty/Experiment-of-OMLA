//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n207), .C1(G1gat), .C2(new_n202), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT17), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(KEYINPUT88), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n214), .A2(KEYINPUT88), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n213), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n216), .B(KEYINPUT15), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n218), .B(new_n219), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n216), .B(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(new_n213), .A3(new_n220), .A4(new_n221), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n219), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n210), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n218), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n209), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n210), .A2(new_n236), .A3(new_n218), .A4(new_n228), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT90), .B1(new_n232), .B2(new_n209), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n231), .B(KEYINPUT13), .Z(new_n240));
  AOI22_X1  g039(.A1(new_n234), .A2(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n233), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n242), .A2(KEYINPUT89), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(KEYINPUT89), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT91), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n242), .B(KEYINPUT89), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n251), .B1(new_n257), .B2(new_n241), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT23), .ZN(new_n267));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(KEYINPUT65), .A3(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n275), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  AND2_X1   g081(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n272), .B(new_n279), .C1(new_n286), .C2(G190gat), .ZN(new_n287));
  AND4_X1   g086(.A1(KEYINPUT25), .A2(new_n265), .A3(new_n267), .A4(new_n268), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n281), .A2(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT67), .A3(new_n263), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(new_n266), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n296), .C1(KEYINPUT26), .C2(new_n263), .ZN(new_n297));
  INV_X1    g096(.A(new_n284), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(KEYINPUT27), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301));
  AOI21_X1  g100(.A(G190gat), .B1(new_n301), .B2(G183gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT28), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n301), .A2(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n297), .B(new_n270), .C1(new_n303), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n263), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n310), .A2(new_n294), .B1(new_n291), .B2(new_n266), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n311), .A2(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n301), .A2(G183gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n277), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n285), .B2(KEYINPUT27), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n316), .B2(KEYINPUT28), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n309), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n290), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G226gat), .ZN(new_n320));
  INV_X1    g119(.A(G233gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n287), .A2(new_n288), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT25), .B1(new_n269), .B2(new_n280), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n322), .B(new_n307), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n328));
  AND2_X1   g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(G211gat), .A2(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G211gat), .ZN(new_n332));
  INV_X1    g131(.A(G218gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  AND4_X1   g142(.A1(new_n331), .A2(new_n337), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n331), .A2(new_n337), .B1(new_n342), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n328), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n337), .A3(new_n342), .A4(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(KEYINPUT76), .A3(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n324), .A2(KEYINPUT77), .A3(new_n327), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n307), .A2(KEYINPUT68), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n317), .A2(new_n309), .A3(new_n270), .A4(new_n297), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n289), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n323), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n327), .B(new_n352), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n361));
  INV_X1    g160(.A(new_n322), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n362), .B(new_n289), .C1(new_n354), .C2(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n357), .B1(new_n290), .B2(new_n307), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n360), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT78), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n360), .A3(new_n365), .ZN(new_n373));
  INV_X1    g172(.A(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n376), .A3(new_n370), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n353), .A2(new_n365), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n360), .A4(new_n368), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n372), .A2(new_n375), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  INV_X1    g180(.A(G120gat), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT69), .B1(new_n382), .B2(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT69), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(G120gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(G113gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT70), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT70), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n383), .A2(new_n386), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  INV_X1    g190(.A(G134gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G127gat), .ZN(new_n393));
  INV_X1    g192(.A(G127gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G134gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n391), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n385), .A2(G120gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n401), .A2(new_n396), .B1(new_n393), .B2(new_n395), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT2), .ZN(new_n406));
  INV_X1    g205(.A(G141gat), .ZN(new_n407));
  INV_X1    g206(.A(G148gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G155gat), .B(G162gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n404), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n397), .B1(new_n388), .B2(KEYINPUT70), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n402), .B1(new_n419), .B2(new_n391), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(new_n412), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n381), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n420), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n415), .B2(new_n416), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n423), .A2(KEYINPUT3), .A3(new_n424), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n404), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n431), .B1(new_n420), .B2(new_n425), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n430), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n381), .B(new_n428), .C1(new_n440), .C2(new_n432), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(KEYINPUT80), .A3(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n430), .B(new_n448), .C1(new_n438), .C2(new_n429), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n449), .ZN(new_n452));
  INV_X1    g251(.A(new_n447), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT6), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n442), .A2(new_n447), .A3(new_n449), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n380), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n356), .A2(new_n404), .ZN(new_n458));
  AOI211_X1 g257(.A(new_n420), .B(new_n289), .C1(new_n354), .C2(new_n355), .ZN(new_n459));
  INV_X1    g258(.A(G227gat), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n458), .A2(new_n459), .B1(new_n460), .B2(new_n321), .ZN(new_n461));
  XOR2_X1   g260(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n460), .A2(new_n321), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT64), .Z(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT34), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n458), .B2(new_n459), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n319), .A2(new_n420), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n356), .A2(new_n404), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT32), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G71gat), .B(G99gat), .Z(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n476), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n482), .B2(new_n480), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(KEYINPUT32), .A3(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n471), .A3(new_n481), .A4(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n461), .A2(new_n465), .A3(new_n462), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n465), .B1(new_n461), .B2(new_n462), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n471), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n481), .A2(new_n485), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g292(.A1(G228gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n349), .A2(new_n496), .A3(new_n350), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n433), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n417), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT3), .B1(new_n423), .B2(new_n424), .ZN(new_n500));
  OAI22_X1  g299(.A1(new_n500), .A2(KEYINPUT29), .B1(new_n344), .B2(new_n345), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n346), .B(new_n351), .C1(new_n500), .C2(KEYINPUT29), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n499), .A3(new_n495), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n498), .B2(new_n417), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT82), .A3(new_n503), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G22gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT84), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(new_n501), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n494), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n507), .A2(KEYINPUT82), .A3(new_n503), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT82), .B1(new_n507), .B2(new_n503), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n510), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT83), .ZN(new_n519));
  OAI21_X1  g318(.A(G22gat), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n511), .B(new_n518), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G50gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n508), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n510), .B1(new_n530), .B2(new_n513), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n493), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT85), .B(new_n532), .C1(new_n523), .C2(new_n526), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n457), .B(new_n492), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n486), .A2(new_n491), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n516), .B(KEYINPUT84), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n509), .A2(new_n519), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(G22gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n528), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT85), .B1(new_n543), .B2(new_n532), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n493), .A3(new_n533), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n380), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n442), .A2(KEYINPUT86), .A3(new_n449), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT86), .B1(new_n442), .B2(new_n449), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n447), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n454), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT35), .B1(new_n551), .B2(new_n450), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n544), .B(new_n545), .C1(new_n456), .C2(new_n380), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n486), .A2(new_n491), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n486), .B2(new_n491), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n438), .A2(new_n429), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n418), .A2(new_n428), .A3(new_n426), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT39), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n453), .C1(KEYINPUT39), .C2(new_n560), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT40), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n380), .A2(new_n550), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n534), .B2(new_n535), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n450), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n289), .B1(new_n317), .B2(new_n312), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n319), .A2(new_n362), .B1(new_n568), .B2(new_n357), .ZN(new_n569));
  INV_X1    g368(.A(new_n327), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n319), .B2(new_n323), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n569), .A2(new_n361), .B1(new_n571), .B2(new_n352), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT38), .B1(new_n572), .B2(KEYINPUT37), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n573), .B(new_n374), .C1(KEYINPUT37), .C2(new_n373), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n374), .A2(KEYINPUT37), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n375), .A2(new_n575), .B1(new_n373), .B2(KEYINPUT37), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT38), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n574), .B(new_n369), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n555), .B(new_n559), .C1(new_n566), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n260), .B1(new_n554), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G57gat), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(G64gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(G64gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(KEYINPUT92), .B2(new_n586), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(KEYINPUT92), .B2(new_n586), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n592), .B1(new_n583), .B2(new_n584), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n593), .A2(new_n597), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n394), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n600), .A2(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n210), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n394), .A3(new_n608), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n610), .B2(new_n614), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  INV_X1    g416(.A(G155gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT96), .B(G92gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(G85gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT8), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G99gat), .B(G106gat), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT7), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n629), .C1(G85gat), .C2(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n632), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n631), .A2(KEYINPUT97), .A3(new_n633), .A4(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n232), .ZN(new_n643));
  NAND3_X1  g442(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n225), .A2(new_n229), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n642), .ZN(new_n646));
  XOR2_X1   g445(.A(G134gat), .B(G162gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G190gat), .B(G218gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT98), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n648), .B(new_n652), .Z(new_n653));
  NAND4_X1  g452(.A1(new_n594), .A2(new_n636), .A3(new_n598), .A4(new_n638), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n611), .B2(new_n642), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n659));
  XOR2_X1   g458(.A(G120gat), .B(G148gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT100), .ZN(new_n661));
  XOR2_X1   g460(.A(G176gat), .B(G204gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT10), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n654), .B(new_n665), .C1(new_n611), .C2(new_n642), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n611), .A2(new_n642), .A3(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n656), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(KEYINPUT99), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n657), .B1(new_n666), .B2(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n658), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT101), .Z(new_n679));
  AOI21_X1  g478(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n625), .A2(new_n653), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n581), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n456), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(G1gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1324gat));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  NAND4_X1  g488(.A1(new_n581), .A2(new_n380), .A3(new_n682), .A4(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G8gat), .B1(new_n683), .B2(new_n547), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n690), .ZN(new_n692));
  MUX2_X1   g491(.A(new_n690), .B(new_n692), .S(KEYINPUT42), .Z(G1325gat));
  OR2_X1    g492(.A1(new_n557), .A2(new_n558), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT105), .ZN(new_n695));
  OAI21_X1  g494(.A(G15gat), .B1(new_n683), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n538), .A2(G15gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n683), .B2(new_n697), .ZN(G1326gat));
  NAND2_X1  g497(.A1(new_n544), .A2(new_n545), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n680), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n625), .A3(new_n653), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n581), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n684), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT45), .Z(new_n707));
  NOR3_X1   g506(.A1(new_n703), .A2(new_n625), .A3(new_n260), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  AOI211_X1 g508(.A(KEYINPUT44), .B(new_n653), .C1(new_n554), .C2(new_n580), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n699), .A2(new_n547), .A3(new_n492), .A4(new_n552), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT35), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n546), .B2(new_n457), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n580), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n653), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n709), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n684), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n722), .ZN(G1328gat));
  OAI21_X1  g522(.A(G36gat), .B1(new_n721), .B2(new_n547), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n705), .A2(G36gat), .A3(new_n547), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(G1329gat));
  NOR3_X1   g526(.A1(new_n705), .A2(G43gat), .A3(new_n538), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n694), .B(new_n708), .C1(new_n710), .C2(new_n718), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n731), .A2(KEYINPUT106), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n695), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n720), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n699), .B1(new_n705), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n741), .B2(new_n705), .ZN(new_n743));
  INV_X1    g542(.A(G50gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n699), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n720), .A2(G50gat), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT48), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1331gat));
  NAND2_X1  g551(.A1(new_n625), .A2(new_n653), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n256), .A2(new_n258), .ZN(new_n754));
  AOI211_X1 g553(.A(KEYINPUT91), .B(new_n251), .C1(new_n257), .C2(new_n241), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n716), .A2(new_n703), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n456), .B(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g560(.A(new_n547), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT109), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT110), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n763), .B(new_n766), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n758), .A2(new_n768), .A3(new_n492), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n758), .A2(new_n737), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n768), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g571(.A1(new_n758), .A2(new_n746), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  INV_X1    g573(.A(new_n625), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n260), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n716), .A2(new_n717), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n680), .A2(new_n684), .A3(G85gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n777), .A2(new_n703), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n710), .B2(new_n718), .ZN(new_n785));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n684), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(G1336gat));
  NOR3_X1   g586(.A1(new_n547), .A2(new_n680), .A3(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n380), .B(new_n784), .C1(new_n710), .C2(new_n718), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n626), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n791), .A2(KEYINPUT111), .A3(new_n626), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT111), .B1(new_n791), .B2(new_n626), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n653), .B(new_n776), .C1(new_n554), .C2(new_n580), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n779), .B1(new_n796), .B2(KEYINPUT112), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n798), .A3(KEYINPUT51), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n797), .A2(new_n799), .A3(new_n788), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n794), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n793), .B1(new_n801), .B2(new_n790), .ZN(G1337gat));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G99gat), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n780), .A2(new_n492), .A3(new_n703), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n785), .A2(new_n695), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n803), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n699), .A2(G106gat), .A3(new_n680), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n780), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n746), .B(new_n784), .C1(new_n710), .C2(new_n718), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(G106gat), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n799), .A3(new_n807), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT115), .B1(new_n816), .B2(KEYINPUT53), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n818), .B(new_n819), .C1(new_n812), .C2(new_n815), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n817), .B2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n674), .A2(new_n822), .A3(new_n676), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n666), .A2(new_n657), .A3(new_n667), .ZN(new_n824));
  AND4_X1   g623(.A1(KEYINPUT117), .A2(new_n669), .A3(KEYINPUT54), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n675), .A2(new_n822), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n826), .B2(new_n824), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n663), .B(new_n823), .C1(new_n825), .C2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n823), .A2(new_n663), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n824), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n826), .A2(KEYINPUT117), .A3(new_n824), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n836), .A3(KEYINPUT55), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n756), .A2(new_n671), .A3(new_n830), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n239), .A2(new_n240), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n231), .B1(new_n230), .B2(new_n233), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n249), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n254), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n703), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n717), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n717), .A2(new_n830), .A3(new_n843), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n671), .B1(new_n828), .B2(new_n829), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n775), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n682), .A2(new_n260), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g650(.A1(new_n547), .A2(new_n851), .A3(new_n546), .A4(new_n759), .ZN(new_n852));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n756), .ZN(new_n853));
  INV_X1    g652(.A(new_n546), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n456), .A3(new_n547), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n385), .A3(new_n260), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n852), .B2(new_n703), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n856), .A2(new_n382), .A3(new_n680), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n852), .A2(new_n394), .A3(new_n625), .ZN(new_n862));
  OAI21_X1  g661(.A(G127gat), .B1(new_n856), .B2(new_n775), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1342gat));
  NAND3_X1  g663(.A1(new_n852), .A2(new_n392), .A3(new_n717), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n856), .B2(new_n653), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  AND2_X1   g668(.A1(new_n851), .A2(new_n759), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n737), .A2(new_n699), .A3(new_n380), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n407), .B1(new_n872), .B2(new_n260), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n694), .A2(new_n684), .A3(new_n380), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n746), .A2(KEYINPUT57), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n845), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(new_n848), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n845), .B2(KEYINPUT118), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n775), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(new_n850), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n699), .B1(new_n849), .B2(new_n850), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n874), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n756), .A2(G141gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n873), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n873), .B(KEYINPUT58), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n408), .A2(KEYINPUT59), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n883), .B2(new_n680), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n699), .A2(KEYINPUT57), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT55), .B1(new_n831), .B2(new_n836), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n847), .A2(new_n894), .A3(new_n260), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n680), .A2(new_n842), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n653), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n625), .B1(new_n897), .B2(new_n877), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n681), .A2(KEYINPUT119), .A3(new_n756), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT119), .B1(new_n681), .B2(new_n756), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n893), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n874), .A2(new_n703), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n902), .B(new_n903), .C1(new_n881), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G148gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n892), .B1(new_n906), .B2(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT120), .B(new_n908), .C1(new_n905), .C2(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n891), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n872), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n408), .A3(new_n703), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n883), .B2(new_n775), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n618), .A3(new_n625), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  INV_X1    g715(.A(G162gat), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n883), .A2(new_n917), .A3(new_n653), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n872), .B2(new_n653), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n547), .A2(new_n456), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n851), .A2(new_n546), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n756), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n759), .A2(new_n547), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n855), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n260), .A2(new_n261), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n922), .A2(new_n262), .A3(new_n703), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n925), .A2(new_n703), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n262), .ZN(G1349gat));
  NAND3_X1  g729(.A1(new_n855), .A2(new_n625), .A3(new_n924), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT121), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n855), .A2(new_n933), .A3(new_n625), .A4(new_n924), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n286), .A3(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n922), .A2(new_n314), .A3(new_n305), .A4(new_n625), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n937), .B(new_n939), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n277), .A3(new_n717), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT123), .Z(new_n942));
  AOI21_X1  g741(.A(new_n277), .B1(new_n925), .B2(new_n717), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n851), .A2(new_n921), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n737), .A2(new_n699), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n756), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n881), .A2(new_n904), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n902), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n695), .A2(new_n924), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n756), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  OAI21_X1  g757(.A(G204gat), .B1(new_n955), .B2(new_n680), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n680), .A2(G204gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n947), .A2(new_n948), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n947), .A2(new_n967), .A3(new_n948), .A4(new_n960), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT125), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n959), .A2(new_n966), .A3(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n332), .A3(new_n625), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n952), .A2(new_n625), .A3(new_n902), .A4(new_n954), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  NAND2_X1  g774(.A1(new_n955), .A2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n952), .A2(new_n977), .A3(new_n902), .A4(new_n954), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(G218gat), .A3(new_n717), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n333), .B1(new_n949), .B2(new_n653), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g781(.A(KEYINPUT126), .B(new_n333), .C1(new_n949), .C2(new_n653), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n976), .A2(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1355gat));
endmodule


