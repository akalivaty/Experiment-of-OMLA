//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT65), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n461), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n465), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n475), .B2(G126), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  NOR2_X1   g067(.A1(KEYINPUT6), .A2(G651), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT6), .A2(G651), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  OAI22_X1  g071(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT66), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n501), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n498), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n495), .A2(new_n496), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n504), .B2(new_n505), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G651), .B1(G50), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n510), .A2(new_n517), .ZN(G166));
  AND3_X1   g093(.A1(new_n498), .A2(G89), .A3(new_n508), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n495), .B2(new_n496), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT67), .B(new_n520), .C1(new_n495), .C2(new_n496), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n528), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n516), .A2(G51), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n519), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(G52), .B2(new_n516), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n498), .A2(G90), .A3(new_n508), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  INV_X1    g114(.A(KEYINPUT68), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n498), .A2(G81), .A3(new_n508), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n516), .A2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n503), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n512), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(G43), .B2(new_n516), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n498), .A2(new_n508), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n549), .B(KEYINPUT68), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n498), .A2(G91), .A3(new_n508), .ZN(new_n560));
  OAI21_X1  g135(.A(G543), .B1(new_n494), .B2(new_n493), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n516), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(KEYINPUT69), .B(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n512), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n560), .A2(new_n566), .A3(new_n570), .ZN(G299));
  OAI21_X1  g146(.A(KEYINPUT70), .B1(new_n519), .B2(new_n531), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n498), .A2(G89), .A3(new_n508), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n573), .A2(new_n574), .A3(new_n525), .A4(new_n530), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n509), .A2(G87), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n501), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n516), .B2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n503), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT71), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(KEYINPUT71), .B1(G48), .B2(new_n516), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n509), .A2(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n503), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT72), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(G47), .B2(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n509), .A2(G85), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n592), .B(new_n593), .C1(new_n591), .C2(new_n590), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT73), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n498), .A2(G92), .A3(new_n508), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n498), .A2(new_n508), .A3(G92), .A4(new_n598), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n516), .A2(G54), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT75), .B(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n512), .A2(new_n604), .B1(new_n605), .B2(new_n515), .ZN(new_n606));
  OAI21_X1  g181(.A(G651), .B1(new_n606), .B2(KEYINPUT76), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n605), .A2(new_n515), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT75), .B(G66), .Z(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n501), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n596), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n596), .B1(G868), .B2(new_n614), .ZN(G321));
  NOR2_X1   g191(.A1(G299), .A2(G868), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n576), .B2(G868), .ZN(G280));
  XNOR2_X1  g193(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n482), .A2(new_n466), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AOI22_X1  g206(.A1(G123), .A2(new_n475), .B1(new_n464), .B2(G135), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n633), .A2(new_n465), .A3(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n465), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n630), .A2(new_n631), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(KEYINPUT80), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(KEYINPUT80), .ZN(new_n647));
  OAI22_X1  g222(.A1(new_n646), .A2(new_n647), .B1(new_n642), .B2(new_n643), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n658), .A2(KEYINPUT81), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(KEYINPUT81), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n629), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n638), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT82), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  INV_X1    g265(.A(new_n688), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n686), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n689), .B2(new_n693), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  AOI22_X1  g273(.A1(G119), .A2(new_n475), .B1(new_n464), .B2(G131), .ZN(new_n699));
  NOR2_X1   g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT83), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G25), .B(new_n703), .S(G29), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n711), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1971), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n711), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT33), .B(G1976), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n710), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n707), .B1(new_n720), .B2(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(G290), .A2(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n711), .A2(G24), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT84), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT85), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1986), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n721), .B(new_n727), .C1(KEYINPUT34), .C2(new_n720), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n482), .A2(G127), .ZN(new_n732));
  AND2_X1   g307(.A1(G115), .A2(G2104), .ZN(new_n733));
  OAI21_X1  g308(.A(G2105), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT25), .ZN(new_n735));
  NAND2_X1  g310(.A1(G103), .A2(G2104), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n464), .A2(G139), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G2072), .Z(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NOR2_X1   g318(.A1(G171), .A2(new_n711), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G5), .B2(new_n711), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n464), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G128), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(new_n748), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2067), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(G2067), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT29), .B(G2090), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n748), .A2(G35), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n479), .B2(G29), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n748), .A2(G32), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n475), .A2(G129), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT26), .Z(new_n769));
  AND3_X1   g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(new_n748), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT89), .ZN(new_n777));
  AOI21_X1  g352(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n637), .B2(new_n748), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n760), .B2(new_n763), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n746), .A2(new_n764), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G160), .A2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n785), .B2(KEYINPUT24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT24), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2084), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT88), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT90), .Z(new_n793));
  NAND3_X1  g368(.A1(new_n783), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n711), .A2(G20), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  INV_X1    g371(.A(G299), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n711), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1956), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n554), .A2(new_n711), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n711), .B2(G19), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n799), .B1(G1341), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G27), .A2(G29), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G164), .B2(G29), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT91), .B(G2078), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n803), .B1(KEYINPUT92), .B2(new_n808), .C1(G1341), .C2(new_n802), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT92), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n711), .A2(G21), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G168), .B2(new_n711), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1966), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n743), .B2(new_n745), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n711), .A2(G4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n614), .B2(new_n711), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G1348), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(G1348), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n810), .A2(new_n814), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n794), .A2(new_n809), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n730), .A2(new_n731), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n499), .B2(new_n500), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(KEYINPUT94), .B(new_n826), .C1(new_n512), .C2(new_n824), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(G651), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n516), .A2(G55), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n498), .A2(G93), .A3(new_n508), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n553), .B2(new_n833), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n614), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n840), .A2(new_n841), .A3(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n844));
  XOR2_X1   g419(.A(new_n843), .B(new_n844), .Z(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(G160), .B(new_n479), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n637), .Z(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n491), .B(new_n755), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n740), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n770), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n703), .B(new_n627), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n475), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n464), .A2(G142), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n856), .A2(new_n465), .A3(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n465), .B2(G118), .ZN(new_n858));
  OR2_X1    g433(.A1(G106), .A2(G2105), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(G2104), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n854), .B(new_n855), .C1(new_n857), .C2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n853), .B(new_n861), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n852), .A2(KEYINPUT97), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(KEYINPUT98), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n852), .A2(new_n862), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(KEYINPUT98), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n849), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n867), .B(new_n849), .C1(new_n862), .C2(new_n852), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(G395));
  INV_X1    g452(.A(G868), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n833), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT99), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n836), .B(new_n622), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n797), .B1(new_n602), .B2(new_n613), .ZN(new_n882));
  INV_X1    g457(.A(new_n603), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n503), .B1(new_n610), .B2(new_n611), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n606), .A2(KEYINPUT76), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n886), .A2(G299), .A3(new_n601), .A4(new_n600), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n888), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n881), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(G166), .B(G288), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n878), .B1(new_n896), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  MUX2_X1   g478(.A(KEYINPUT99), .B(new_n880), .S(new_n903), .Z(G295));
  MUX2_X1   g479(.A(KEYINPUT99), .B(new_n880), .S(new_n903), .Z(G331));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n572), .A2(G171), .A3(new_n575), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(G168), .B2(G301), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n572), .A2(G171), .A3(new_n908), .A4(new_n575), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n836), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n553), .A2(new_n833), .ZN(new_n913));
  INV_X1    g488(.A(new_n835), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n910), .A2(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n892), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT101), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n892), .B(new_n918), .C1(new_n912), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n912), .A2(new_n894), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n572), .A2(G171), .A3(new_n575), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n573), .A2(new_n525), .A3(new_n530), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT100), .B1(G171), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n911), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n913), .A2(new_n914), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n915), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n900), .B1(new_n920), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n906), .B1(new_n932), .B2(G37), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n928), .A2(new_n930), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n917), .A2(new_n919), .B1(new_n934), .B2(new_n921), .ZN(new_n935));
  OAI211_X1 g510(.A(KEYINPUT103), .B(new_n873), .C1(new_n935), .C2(new_n900), .ZN(new_n936));
  INV_X1    g511(.A(new_n919), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n836), .A2(new_n910), .A3(new_n911), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n918), .B1(new_n939), .B2(new_n892), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n931), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT104), .B1(new_n941), .B2(new_n899), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n920), .A2(new_n943), .A3(new_n900), .A4(new_n931), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n933), .A2(new_n936), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n899), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT103), .B1(new_n949), .B2(new_n873), .ZN(new_n950));
  AOI211_X1 g525(.A(new_n906), .B(G37), .C1(new_n941), .C2(new_n899), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n921), .A2(new_n927), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n928), .A2(new_n938), .A3(new_n930), .ZN(new_n957));
  INV_X1    g532(.A(new_n892), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n899), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n948), .A2(new_n960), .A3(new_n946), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n947), .A2(new_n954), .A3(new_n955), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n948), .A2(new_n946), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n936), .B2(new_n933), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n946), .B1(new_n948), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n962), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n491), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G1996), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT46), .Z(new_n974));
  XOR2_X1   g549(.A(new_n972), .B(KEYINPUT106), .Z(new_n975));
  XNOR2_X1  g550(.A(new_n755), .B(G2067), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n770), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n982), .B2(new_n770), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n983), .A2(new_n975), .B1(new_n770), .B2(new_n973), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n703), .A2(new_n706), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n703), .A2(new_n706), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n972), .A2(G1986), .A3(G290), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n981), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(new_n985), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G2067), .B2(new_n755), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n975), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT63), .ZN(new_n995));
  OAI211_X1 g570(.A(G303), .B(G8), .C1(KEYINPUT109), .C2(KEYINPUT55), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(G166), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n491), .A2(new_n968), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n970), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n969), .A2(new_n970), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1971), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(G8), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1000), .B(G8), .C1(new_n1009), .C2(new_n1006), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n971), .A2(new_n968), .A3(new_n491), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT110), .B1(G288), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n579), .A2(new_n1026), .A3(G1976), .A4(new_n581), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1025), .A2(new_n1014), .A3(G8), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1032), .A3(KEYINPUT52), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1028), .B2(KEYINPUT52), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1023), .B(new_n1031), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1013), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(G2084), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1042));
  INV_X1    g617(.A(G1966), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1003), .A2(new_n1005), .A3(KEYINPUT114), .A4(new_n789), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G286), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n995), .B1(new_n1038), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT63), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1036), .A2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1021), .A2(new_n1022), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(KEYINPUT112), .C1(new_n1035), .C2(new_n1034), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1056), .A2(KEYINPUT115), .A3(new_n1048), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n1056), .B2(new_n1048), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1050), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1012), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1060));
  XOR2_X1   g635(.A(new_n1015), .B(KEYINPUT113), .Z(new_n1061));
  NAND3_X1  g636(.A1(new_n1023), .A2(new_n1024), .A3(new_n716), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1018), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1046), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1041), .A2(new_n1044), .A3(KEYINPUT123), .A4(new_n1045), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G168), .A2(new_n997), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(G168), .A3(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n997), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1047), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1066), .B(new_n1072), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1073), .A2(new_n1077), .B1(new_n1047), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1072), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT62), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1007), .A2(new_n1085), .A3(new_n1008), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1087), .A2(KEYINPUT53), .B1(new_n743), .B2(new_n1040), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT126), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT126), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1081), .A2(new_n1084), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1956), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1040), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n969), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n1008), .A3(new_n971), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1007), .A2(KEYINPUT119), .A3(new_n1008), .A4(new_n1101), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n560), .A2(new_n570), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1107), .A2(KEYINPUT116), .B1(new_n563), .B2(new_n565), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n560), .A2(new_n1109), .A3(new_n570), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1111), .A2(new_n1112), .B1(KEYINPUT57), .B2(new_n797), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(KEYINPUT120), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n797), .A2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1125), .B2(new_n1116), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1106), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1099), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1130), .A2(G1348), .B1(G2067), .B2(new_n1014), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n614), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1125), .A2(new_n1106), .A3(new_n1116), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT121), .B(KEYINPUT61), .C1(new_n1129), .C2(new_n1135), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(G1348), .ZN(new_n1141));
  INV_X1    g716(.A(G2067), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1014), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1040), .A2(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n614), .A2(KEYINPUT122), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n614), .A2(KEYINPUT122), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1144), .A2(KEYINPUT60), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1147), .B(new_n1149), .C1(new_n1150), .C2(new_n1145), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT58), .B(G1341), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1042), .A2(G1996), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n554), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1153), .A2(new_n1156), .A3(new_n554), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1129), .A2(KEYINPUT61), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1127), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1133), .B1(new_n1140), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1088), .B(G301), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1095), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1094), .B2(G171), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1095), .A2(new_n1163), .A3(new_n1166), .A4(KEYINPUT54), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1168), .B(new_n1169), .C1(new_n1083), .C2(new_n1082), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1097), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1038), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1065), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(G290), .B(G1986), .Z(new_n1174));
  OAI211_X1 g749(.A(new_n984), .B(new_n987), .C1(new_n972), .C2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT108), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n994), .B1(new_n1173), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g752(.A1(G227), .A2(new_n459), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n695), .B2(new_n696), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1180), .A2(G401), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1181), .B1(new_n871), .B2(new_n874), .ZN(new_n1182));
  INV_X1    g756(.A(new_n961), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n1184), .B2(KEYINPUT105), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1185), .B2(new_n954), .ZN(G308));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n954), .ZN(new_n1187));
  INV_X1    g761(.A(new_n1182), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1188), .ZN(G225));
endmodule


