//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1020,
    new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(KEYINPUT66), .A2(KEYINPUT26), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT26), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n217), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n221), .A2(new_n217), .A3(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT28), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n215), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n205), .A2(new_n233), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n206), .A2(new_n210), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(KEYINPUT24), .A3(new_n204), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT25), .A4(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n234), .A2(new_n231), .A3(new_n230), .A4(new_n236), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n215), .A2(new_n226), .A3(new_n242), .A4(new_n227), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n229), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G127gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G134gat), .ZN(new_n246));
  INV_X1    g045(.A(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G127gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT68), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(new_n247), .A3(G127gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(new_n245), .B2(G134gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n247), .A2(G127gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n253), .A4(new_n259), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n256), .A2(new_n258), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n271));
  OR3_X1    g070(.A1(new_n257), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n246), .A2(new_n248), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n274));
  AND4_X1   g073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n203), .B1(new_n244), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n228), .A2(KEYINPUT67), .B1(new_n240), .B2(new_n237), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n262), .B2(new_n268), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT73), .A4(new_n243), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n244), .A2(new_n277), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT74), .B(KEYINPUT33), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT75), .ZN(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  NAND3_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n278), .A2(new_n284), .A3(new_n281), .A4(new_n282), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT34), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT34), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(new_n283), .B2(new_n285), .ZN(new_n301));
  INV_X1    g100(.A(new_n288), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n283), .B2(new_n285), .ZN(new_n303));
  INV_X1    g102(.A(new_n293), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n294), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT78), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT78), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n294), .A2(new_n299), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n311));
  AOI221_X4 g110(.A(new_n300), .B1(new_n302), .B2(new_n293), .C1(new_n283), .C2(new_n285), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT76), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n299), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n315), .A3(new_n305), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n202), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n299), .B1(new_n294), .B2(new_n305), .ZN(new_n319));
  AOI211_X1 g118(.A(KEYINPUT36), .B(new_n319), .C1(new_n307), .C2(new_n309), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n244), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327));
  OR2_X1    g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  NAND2_X1  g129(.A1(G211gat), .A2(G218gat), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n332), .B2(new_n333), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n327), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n328), .A2(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n330), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT79), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(KEYINPUT80), .A3(new_n334), .A4(new_n337), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n342), .B2(new_n337), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n332), .A2(KEYINPUT81), .A3(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n325), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n244), .B2(new_n322), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n241), .A2(new_n228), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n351), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT82), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n326), .B(new_n350), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n322), .A3(new_n325), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n244), .B2(new_n325), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n349), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  AND3_X1   g161(.A1(new_n356), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n356), .B2(new_n359), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n356), .A2(new_n359), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n367), .A2(new_n365), .A3(new_n362), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  XOR2_X1   g169(.A(G141gat), .B(G148gat), .Z(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT2), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n372), .B1(new_n371), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT83), .A3(new_n376), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT3), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT84), .A4(KEYINPUT3), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n377), .A2(new_n378), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n277), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n280), .B2(new_n386), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n280), .A2(new_n391), .A3(new_n386), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n389), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n390), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n381), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n280), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n376), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n275), .B(new_n398), .C1(new_n262), .C2(new_n268), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n399), .A2(new_n391), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n280), .A2(new_n386), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n390), .A4(new_n389), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n402), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT92), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n412), .A3(new_n415), .A4(new_n407), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(KEYINPUT91), .A2(KEYINPUT40), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT90), .B(KEYINPUT39), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n395), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n390), .B1(new_n411), .B2(new_n389), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n280), .B2(new_n396), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT39), .B1(new_n423), .B2(new_n395), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(new_n406), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(KEYINPUT91), .A2(KEYINPUT40), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n369), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT86), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n346), .A2(new_n433), .A3(new_n347), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n342), .A2(new_n337), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n346), .B2(new_n347), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n322), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n386), .B1(new_n438), .B2(new_n387), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n386), .B2(new_n387), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n349), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n349), .A2(new_n322), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n396), .B1(new_n443), .B2(new_n387), .ZN(new_n444));
  OAI211_X1 g243(.A(G228gat), .B(G233gat), .C1(new_n349), .C2(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT88), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n388), .A2(new_n322), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n431), .B1(new_n350), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n349), .B2(new_n322), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n448), .B(new_n449), .C1(new_n396), .C2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G22gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n452), .A2(new_n455), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n457), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n456), .B2(new_n457), .ZN(new_n464));
  AOI211_X1 g263(.A(KEYINPUT89), .B(G22gat), .C1(new_n452), .C2(new_n455), .ZN(new_n465));
  OAI22_X1  g264(.A1(new_n464), .A2(new_n465), .B1(new_n452), .B2(new_n455), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n356), .A2(new_n468), .A3(new_n359), .ZN(new_n469));
  INV_X1    g268(.A(new_n362), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n326), .B(new_n349), .C1(new_n352), .C2(new_n355), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n358), .B2(new_n350), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT38), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n363), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n367), .A2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n470), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n413), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n402), .A2(new_n412), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n406), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n414), .A2(new_n482), .A3(new_n479), .A4(new_n416), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n475), .A2(new_n478), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n430), .A2(new_n467), .A3(new_n484), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n367), .A2(new_n365), .A3(new_n362), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n482), .A2(new_n489), .A3(new_n479), .A4(new_n413), .ZN(new_n490));
  INV_X1    g289(.A(new_n481), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(new_n407), .C1(KEYINPUT85), .C2(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n466), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n321), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n319), .B1(new_n307), .B2(new_n309), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n467), .A2(new_n499), .A3(new_n488), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT35), .B1(new_n483), .B2(new_n480), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n487), .A2(new_n486), .B1(new_n490), .B2(new_n492), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n467), .A2(new_n502), .A3(new_n310), .A4(new_n317), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n500), .A2(new_n501), .B1(new_n503), .B2(KEYINPUT35), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G197gat), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT11), .B(G169gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT12), .Z(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT13), .Z(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n461), .A2(G15gat), .ZN(new_n514));
  INV_X1    g313(.A(G15gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G22gat), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT94), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT94), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(G1gat), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n515), .A2(G22gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n461), .A2(G15gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT94), .ZN(new_n526));
  AOI21_X1  g325(.A(G1gat), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(KEYINPUT95), .B(new_n513), .C1(new_n521), .C2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n525), .B(new_n526), .C1(new_n519), .C2(G1gat), .ZN(new_n529));
  INV_X1    g328(.A(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n517), .B2(new_n518), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n513), .A2(KEYINPUT95), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n513), .A2(KEYINPUT95), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n536), .B2(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(G29gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT15), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(new_n537), .C1(new_n539), .C2(new_n541), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n549), .A3(KEYINPUT15), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n547), .B2(new_n550), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n535), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT93), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n555), .A2(new_n556), .B1(new_n528), .B2(new_n534), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n512), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n528), .A4(new_n534), .ZN(new_n559));
  NOR3_X1   g358(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT17), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n547), .A2(KEYINPUT17), .A3(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n511), .B(new_n559), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT18), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n555), .A2(new_n566), .A3(new_n556), .ZN(new_n567));
  INV_X1    g366(.A(new_n550), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n549), .B1(new_n542), .B2(KEYINPUT15), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n545), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n570), .A2(KEYINPUT17), .B1(new_n528), .B2(new_n534), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n551), .A2(new_n552), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n528), .A2(new_n534), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n567), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT18), .B1(new_n574), .B2(new_n511), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n510), .B1(new_n565), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(KEYINPUT18), .A3(new_n511), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n563), .A2(new_n564), .ZN(new_n578));
  INV_X1    g377(.A(new_n510), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n558), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT97), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n586), .B2(KEYINPUT9), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT97), .ZN(new_n589));
  INV_X1    g388(.A(G57gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(G64gat), .ZN(new_n591));
  INV_X1    g390(.A(G64gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G57gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(KEYINPUT96), .A2(G71gat), .A3(G78gat), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n597), .A2(new_n598), .A3(new_n586), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n588), .B(new_n584), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n591), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n592), .A2(G57gat), .ZN(new_n604));
  OR2_X1    g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(KEYINPUT98), .A2(new_n604), .B1(new_n605), .B2(new_n585), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n535), .B1(new_n583), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT99), .B(KEYINPUT19), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n583), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT20), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(new_n614), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G183gat), .B(G211gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n624), .B1(new_n619), .B2(new_n622), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n612), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n611), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G99gat), .B(G106gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT7), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(KEYINPUT100), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT8), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n634), .B1(new_n639), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT7), .ZN(new_n649));
  AOI22_X1  g448(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n649), .A2(new_n633), .A3(new_n641), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n567), .A2(new_n561), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n648), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n555), .A2(new_n556), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n656));
  INV_X1    g455(.A(G232gat), .ZN(new_n657));
  INV_X1    g456(.A(G233gat), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(KEYINPUT101), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT101), .B1(new_n655), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n653), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G190gat), .B(G218gat), .Z(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n655), .A2(new_n660), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n661), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n667), .B1(new_n671), .B2(new_n653), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI22_X1  g476(.A1(new_n666), .A2(new_n672), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n664), .A2(new_n665), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n671), .A2(new_n667), .A3(new_n653), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n677), .A2(new_n673), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n651), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n607), .A3(new_n600), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n654), .ZN(new_n687));
  INV_X1    g486(.A(G230gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n658), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n605), .A2(new_n585), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n604), .A2(KEYINPUT98), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n603), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n692), .A2(new_n601), .B1(new_n595), .B2(new_n599), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n652), .A3(new_n685), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n687), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n696));
  INV_X1    g495(.A(new_n689), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT10), .B1(new_n687), .B2(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT10), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n608), .A2(new_n652), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(G120gat), .B(G148gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(G176gat), .B(G204gat), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n695), .A2(KEYINPUT104), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n696), .A2(new_n701), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n701), .B2(new_n695), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n632), .A2(new_n678), .A3(new_n683), .A4(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n505), .A2(new_n582), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n493), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g513(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n519), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(new_n369), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n717), .A2(G8gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(G8gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n711), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n488), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n718), .B(new_n719), .C1(KEYINPUT42), .C2(new_n721), .ZN(G1325gat));
  NOR2_X1   g521(.A1(new_n318), .A2(new_n320), .ZN(new_n723));
  OAI21_X1  g522(.A(G15gat), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n711), .A2(new_n515), .A3(new_n499), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n495), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  NOR2_X1   g528(.A1(new_n505), .A2(new_n582), .ZN(new_n730));
  INV_X1    g529(.A(new_n709), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n632), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n678), .A2(new_n683), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n730), .A2(new_n536), .A3(new_n712), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT45), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n734), .A2(KEYINPUT44), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n498), .B2(new_n504), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n576), .A2(KEYINPUT106), .A3(new_n580), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT106), .B1(new_n576), .B2(new_n580), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n496), .A2(KEYINPUT107), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n494), .A2(new_n495), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n723), .A2(new_n745), .A3(new_n485), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n467), .A2(new_n499), .A3(new_n488), .A4(new_n501), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n735), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n740), .B(new_n744), .C1(new_n752), .C2(KEYINPUT44), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(KEYINPUT108), .A3(new_n493), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n753), .B2(new_n493), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G29gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n738), .B1(new_n754), .B2(new_n756), .ZN(G1328gat));
  NAND4_X1  g556(.A1(new_n730), .A2(new_n538), .A3(new_n369), .A4(new_n736), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g558(.A(G36gat), .B1(new_n753), .B2(new_n488), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(G1329gat));
  OAI21_X1  g561(.A(G43gat), .B1(new_n753), .B2(new_n723), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  INV_X1    g563(.A(new_n499), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(G43gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n730), .A2(new_n736), .A3(new_n766), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(new_n763), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1330gat));
  OAI21_X1  g569(.A(G50gat), .B1(new_n753), .B2(new_n467), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n467), .A2(G50gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n730), .A2(new_n736), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n771), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(G1331gat));
  NAND2_X1  g576(.A1(new_n748), .A2(new_n751), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n581), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n576), .A2(KEYINPUT106), .A3(new_n580), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n632), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n782), .A2(new_n734), .A3(new_n783), .A4(new_n709), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n493), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(new_n590), .ZN(G1332gat));
  AND3_X1   g586(.A1(new_n778), .A2(KEYINPUT109), .A3(new_n784), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT109), .B1(new_n778), .B2(new_n784), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n369), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT49), .B(G64gat), .Z(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(G1333gat));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795));
  INV_X1    g594(.A(G71gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n790), .B2(new_n321), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n785), .A2(G71gat), .A3(new_n765), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n499), .A2(new_n796), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n788), .A2(new_n789), .A3(new_n723), .ZN(new_n801));
  OAI221_X1 g600(.A(KEYINPUT50), .B1(new_n785), .B2(new_n800), .C1(new_n801), .C2(new_n796), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(G1334gat));
  NAND2_X1  g602(.A1(new_n790), .A2(new_n495), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g604(.A1(new_n743), .A2(new_n783), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT110), .ZN(new_n807));
  AND4_X1   g606(.A1(KEYINPUT51), .A2(new_n778), .A3(new_n734), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n752), .B2(new_n807), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n642), .A3(new_n712), .A4(new_n731), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n807), .A2(new_n731), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n740), .B(new_n812), .C1(new_n752), .C2(KEYINPUT44), .ZN(new_n813));
  OAI21_X1  g612(.A(G85gat), .B1(new_n813), .B2(new_n493), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(G1336gat));
  OAI21_X1  g614(.A(G92gat), .B1(new_n813), .B2(new_n488), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n369), .A2(new_n643), .A3(new_n731), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT112), .Z(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n808), .B2(new_n809), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT52), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n816), .B(new_n819), .C1(new_n821), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1337gat));
  NOR3_X1   g625(.A1(new_n765), .A2(G99gat), .A3(new_n709), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G99gat), .B1(new_n813), .B2(new_n723), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1338gat));
  OAI21_X1  g629(.A(G106gat), .B1(new_n813), .B2(new_n467), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n467), .A2(G106gat), .A3(new_n709), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n808), .B2(new_n809), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT113), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  AND4_X1   g637(.A1(new_n632), .A2(new_n678), .A3(new_n683), .A4(new_n709), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT114), .A3(new_n743), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n782), .B2(new_n710), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n686), .A2(new_n654), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n652), .B1(new_n693), .B2(new_n685), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n699), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n700), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n689), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n701), .A3(KEYINPUT54), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n697), .C1(new_n698), .C2(new_n700), .ZN(new_n851));
  INV_X1    g650(.A(new_n704), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT55), .B(new_n849), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n706), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n852), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT55), .B1(new_n861), .B2(new_n849), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n574), .A2(new_n511), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n553), .A2(new_n557), .A3(new_n512), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n509), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n580), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n734), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n731), .A2(new_n867), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n863), .B2(new_n782), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n870), .B2(new_n734), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n843), .B1(new_n871), .B2(new_n783), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n493), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n310), .A2(new_n317), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n467), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n488), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT116), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n257), .A3(new_n782), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n500), .ZN(new_n879));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n582), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1340gat));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n255), .A3(new_n731), .ZN(new_n882));
  OAI21_X1  g681(.A(G120gat), .B1(new_n879), .B2(new_n709), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1341gat));
  OAI21_X1  g683(.A(G127gat), .B1(new_n879), .B2(new_n783), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n632), .A2(new_n245), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n876), .B2(new_n886), .ZN(G1342gat));
  OR3_X1    g686(.A1(new_n876), .A2(G134gat), .A3(new_n735), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n879), .B2(new_n735), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n723), .A2(new_n495), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT120), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n488), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n582), .A2(G141gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n848), .A2(new_n701), .A3(KEYINPUT54), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n859), .B2(new_n860), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n707), .B1(new_n900), .B2(KEYINPUT55), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT55), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n901), .B(new_n904), .C1(new_n741), .C2(new_n742), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n731), .A2(new_n867), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n734), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n863), .A2(new_n734), .A3(new_n867), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n783), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n840), .A2(new_n842), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n467), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n902), .A2(new_n914), .A3(new_n903), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n902), .B2(new_n903), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n582), .A2(new_n856), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n869), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n868), .B1(new_n919), .B2(new_n734), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n843), .B1(new_n920), .B2(new_n783), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n495), .A2(KEYINPUT57), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n911), .A2(new_n913), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n723), .A2(new_n712), .A3(new_n488), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n581), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G141gat), .ZN(new_n927));
  XOR2_X1   g726(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n928));
  NAND3_X1  g727(.A1(new_n898), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n923), .B2(new_n925), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n930), .A3(new_n925), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n782), .A3(new_n933), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n934), .A2(G141gat), .B1(new_n896), .B2(new_n897), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(G1344gat));
  INV_X1    g736(.A(G148gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n896), .A2(new_n938), .A3(new_n731), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n912), .B1(new_n872), .B2(new_n467), .ZN(new_n940));
  INV_X1    g739(.A(new_n922), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n902), .A2(new_n914), .A3(new_n903), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n581), .A3(new_n901), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n906), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n735), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n632), .B1(new_n946), .B2(new_n868), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n947), .B2(new_n843), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT119), .B(new_n924), .C1(new_n940), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n931), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT59), .B(new_n938), .C1(new_n950), .C2(new_n731), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n920), .A2(new_n783), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n581), .B2(new_n710), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n495), .ZN(new_n955));
  INV_X1    g754(.A(new_n911), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n955), .A2(KEYINPUT57), .B1(new_n956), .B2(new_n912), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n731), .A3(new_n925), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n952), .B1(new_n958), .B2(G148gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n939), .B1(new_n951), .B2(new_n959), .ZN(G1345gat));
  AOI21_X1  g759(.A(G155gat), .B1(new_n896), .B2(new_n632), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n632), .A2(G155gat), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT122), .Z(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n950), .B2(new_n963), .ZN(G1346gat));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n374), .B1(new_n950), .B2(new_n734), .ZN(new_n966));
  NOR4_X1   g765(.A1(new_n894), .A2(new_n895), .A3(G162gat), .A4(new_n735), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n896), .A2(new_n374), .A3(new_n734), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n949), .A2(new_n931), .A3(new_n735), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n969), .B(KEYINPUT123), .C1(new_n970), .C2(new_n374), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1347gat));
  NOR2_X1   g771(.A1(new_n712), .A2(new_n488), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n872), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n975), .A2(new_n875), .ZN(new_n976));
  AOI21_X1  g775(.A(G169gat), .B1(new_n976), .B2(new_n782), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(new_n467), .A3(new_n499), .ZN(new_n978));
  INV_X1    g777(.A(G169gat), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(new_n582), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n977), .A2(new_n980), .ZN(G1348gat));
  INV_X1    g780(.A(G176gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n976), .A2(new_n982), .A3(new_n731), .ZN(new_n983));
  OAI21_X1  g782(.A(G176gat), .B1(new_n978), .B2(new_n709), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1349gat));
  NAND4_X1  g784(.A1(new_n976), .A2(new_n207), .A3(new_n209), .A4(new_n632), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n987), .B1(new_n978), .B2(new_n783), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G183gat), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n978), .A2(new_n987), .A3(new_n783), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g791(.A(new_n210), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n978), .B2(new_n735), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI221_X1 g795(.A(new_n993), .B1(KEYINPUT125), .B2(KEYINPUT61), .C1(new_n978), .C2(new_n735), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n976), .A2(new_n210), .A3(new_n734), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g799(.A1(new_n723), .A2(new_n973), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n957), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(G197gat), .ZN(new_n1004));
  NOR3_X1   g803(.A1(new_n1003), .A2(new_n1004), .A3(new_n582), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n956), .A2(new_n1001), .ZN(new_n1006));
  AOI21_X1  g805(.A(G197gat), .B1(new_n1006), .B2(new_n782), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1005), .A2(new_n1007), .ZN(G1352gat));
  XOR2_X1   g807(.A(KEYINPUT127), .B(G204gat), .Z(new_n1009));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n731), .A3(new_n1009), .ZN(new_n1010));
  XOR2_X1   g809(.A(new_n1010), .B(KEYINPUT62), .Z(new_n1011));
  AND3_X1   g810(.A1(new_n957), .A2(new_n731), .A3(new_n1002), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n1012), .B2(new_n1009), .ZN(G1353gat));
  INV_X1    g812(.A(G211gat), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1006), .A2(new_n1014), .A3(new_n632), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n957), .A2(new_n632), .A3(new_n1002), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1016), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1016), .B2(G211gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(G1354gat));
  OAI21_X1  g818(.A(G218gat), .B1(new_n1003), .B2(new_n735), .ZN(new_n1020));
  INV_X1    g819(.A(G218gat), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n1021), .A3(new_n734), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1020), .A2(new_n1022), .ZN(G1355gat));
endmodule


