

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762;

  NOR2_X1 U380 ( .A1(n540), .A2(n379), .ZN(n512) );
  INV_X4 U381 ( .A(G953), .ZN(n752) );
  XNOR2_X1 U382 ( .A(n388), .B(n369), .ZN(n761) );
  XOR2_X1 U383 ( .A(n365), .B(n489), .Z(n357) );
  AND2_X2 U384 ( .A1(n375), .A2(n542), .ZN(n543) );
  AND2_X2 U385 ( .A1(n406), .A2(n410), .ZN(n375) );
  NAND2_X2 U386 ( .A1(n397), .A2(n380), .ZN(n396) );
  AND2_X2 U387 ( .A1(n391), .A2(n761), .ZN(n527) );
  XNOR2_X2 U388 ( .A(KEYINPUT71), .B(G131), .ZN(n457) );
  XNOR2_X2 U389 ( .A(n447), .B(KEYINPUT4), .ZN(n387) );
  INV_X1 U390 ( .A(n611), .ZN(n692) );
  INV_X4 U391 ( .A(G104), .ZN(n403) );
  NAND2_X1 U392 ( .A1(n377), .A2(n367), .ZN(n668) );
  XNOR2_X1 U393 ( .A(n371), .B(KEYINPUT36), .ZN(n558) );
  NAND2_X1 U394 ( .A1(n583), .A2(n485), .ZN(n405) );
  XNOR2_X1 U395 ( .A(n399), .B(n385), .ZN(n611) );
  XNOR2_X1 U396 ( .A(n498), .B(n750), .ZN(n733) );
  INV_X1 U397 ( .A(n377), .ZN(n358) );
  NAND2_X1 U398 ( .A1(n619), .A2(n362), .ZN(n359) );
  AND2_X1 U399 ( .A1(n359), .A2(n360), .ZN(n625) );
  OR2_X1 U400 ( .A1(n361), .A2(n621), .ZN(n360) );
  INV_X1 U401 ( .A(n624), .ZN(n361) );
  AND2_X1 U402 ( .A1(n664), .A2(n624), .ZN(n362) );
  OR2_X1 U403 ( .A1(n557), .A2(n556), .ZN(n371) );
  XNOR2_X1 U404 ( .A(n454), .B(KEYINPUT10), .ZN(n497) );
  XNOR2_X1 U405 ( .A(G146), .B(G125), .ZN(n454) );
  NAND2_X1 U406 ( .A1(n417), .A2(n570), .ZN(n416) );
  INV_X1 U407 ( .A(n677), .ZN(n417) );
  INV_X1 U408 ( .A(G902), .ZN(n510) );
  OR2_X1 U409 ( .A1(n634), .A2(G902), .ZN(n384) );
  XOR2_X1 U410 ( .A(G137), .B(G140), .Z(n505) );
  NAND2_X1 U411 ( .A1(n675), .A2(n674), .ZN(n671) );
  NOR2_X1 U412 ( .A1(n733), .A2(G902), .ZN(n414) );
  XNOR2_X1 U413 ( .A(n422), .B(G107), .ZN(n470) );
  INV_X1 U414 ( .A(G116), .ZN(n422) );
  XNOR2_X1 U415 ( .A(KEYINPUT78), .B(KEYINPUT94), .ZN(n489) );
  XNOR2_X1 U416 ( .A(n423), .B(G110), .ZN(n493) );
  INV_X1 U417 ( .A(G119), .ZN(n423) );
  XNOR2_X1 U418 ( .A(KEYINPUT85), .B(KEYINPUT93), .ZN(n492) );
  XNOR2_X1 U419 ( .A(G128), .B(KEYINPUT24), .ZN(n491) );
  XNOR2_X1 U420 ( .A(n413), .B(n411), .ZN(n488) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n413) );
  NOR2_X1 U422 ( .A1(n412), .A2(G953), .ZN(n411) );
  INV_X1 U423 ( .A(G234), .ZN(n412) );
  XNOR2_X1 U424 ( .A(n497), .B(n456), .ZN(n460) );
  XNOR2_X1 U425 ( .A(n430), .B(n458), .ZN(n459) );
  XOR2_X1 U426 ( .A(G113), .B(G143), .Z(n430) );
  AND2_X1 U427 ( .A1(n644), .A2(n552), .ZN(n555) );
  INV_X1 U428 ( .A(n574), .ZN(n393) );
  INV_X1 U429 ( .A(n692), .ZN(n390) );
  XNOR2_X1 U430 ( .A(n466), .B(n373), .ZN(n570) );
  XNOR2_X1 U431 ( .A(n374), .B(KEYINPUT13), .ZN(n373) );
  INV_X1 U432 ( .A(G475), .ZN(n374) );
  INV_X1 U433 ( .A(KEYINPUT1), .ZN(n385) );
  BUF_X1 U434 ( .A(n686), .Z(n379) );
  INV_X1 U435 ( .A(KEYINPUT103), .ZN(n408) );
  NOR2_X1 U436 ( .A1(n643), .A2(n366), .ZN(n410) );
  INV_X1 U437 ( .A(KEYINPUT73), .ZN(n400) );
  XNOR2_X1 U438 ( .A(G119), .B(G116), .ZN(n434) );
  XNOR2_X1 U439 ( .A(KEYINPUT5), .B(G137), .ZN(n433) );
  XNOR2_X1 U440 ( .A(n457), .B(G134), .ZN(n383) );
  XNOR2_X1 U441 ( .A(G902), .B(KEYINPUT91), .ZN(n441) );
  XNOR2_X1 U442 ( .A(G101), .B(G110), .ZN(n502) );
  XOR2_X1 U443 ( .A(G104), .B(G107), .Z(n503) );
  XNOR2_X1 U444 ( .A(n472), .B(n395), .ZN(n394) );
  XNOR2_X1 U445 ( .A(G146), .B(G125), .ZN(n395) );
  XOR2_X1 U446 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n474) );
  NOR2_X1 U447 ( .A1(n751), .A2(KEYINPUT2), .ZN(n419) );
  INV_X1 U448 ( .A(KEYINPUT86), .ZN(n418) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n480) );
  XNOR2_X1 U450 ( .A(n614), .B(n376), .ZN(n569) );
  INV_X1 U451 ( .A(KEYINPUT38), .ZN(n376) );
  NAND2_X1 U452 ( .A1(n686), .A2(n687), .ZN(n693) );
  XNOR2_X1 U453 ( .A(n401), .B(G101), .ZN(n471) );
  XNOR2_X1 U454 ( .A(KEYINPUT3), .B(G113), .ZN(n401) );
  XNOR2_X1 U455 ( .A(G134), .B(G122), .ZN(n445) );
  XNOR2_X1 U456 ( .A(KEYINPUT9), .B(KEYINPUT101), .ZN(n382) );
  NOR2_X1 U457 ( .A1(n578), .A2(n399), .ZN(n584) );
  NOR2_X1 U458 ( .A1(n671), .A2(n416), .ZN(n573) );
  INV_X1 U459 ( .A(KEYINPUT0), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n424), .B(n421), .ZN(n739) );
  XOR2_X1 U461 ( .A(n493), .B(n470), .Z(n421) );
  XNOR2_X1 U462 ( .A(n402), .B(n471), .ZN(n424) );
  XNOR2_X1 U463 ( .A(n469), .B(KEYINPUT16), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n490), .B(n357), .ZN(n496) );
  XNOR2_X1 U465 ( .A(n363), .B(n463), .ZN(n464) );
  XNOR2_X1 U466 ( .A(n460), .B(n459), .ZN(n465) );
  NOR2_X1 U467 ( .A1(n752), .A2(G952), .ZN(n737) );
  XNOR2_X1 U468 ( .A(n427), .B(n425), .ZN(n762) );
  XNOR2_X1 U469 ( .A(n426), .B(KEYINPUT109), .ZN(n425) );
  AND2_X1 U470 ( .A1(n703), .A2(n584), .ZN(n427) );
  INV_X1 U471 ( .A(KEYINPUT42), .ZN(n426) );
  BUF_X1 U472 ( .A(n525), .Z(n642) );
  AND2_X1 U473 ( .A1(n553), .A2(n390), .ZN(n389) );
  AND2_X1 U474 ( .A1(n512), .A2(n392), .ZN(n641) );
  XOR2_X1 U475 ( .A(n462), .B(n461), .Z(n363) );
  XNOR2_X1 U476 ( .A(KEYINPUT25), .B(KEYINPUT95), .ZN(n364) );
  XOR2_X1 U477 ( .A(KEYINPUT72), .B(KEYINPUT23), .Z(n365) );
  AND2_X1 U478 ( .A1(n672), .A2(KEYINPUT103), .ZN(n366) );
  AND2_X1 U479 ( .A1(n751), .A2(KEYINPUT2), .ZN(n367) );
  NOR2_X1 U480 ( .A1(n672), .A2(KEYINPUT103), .ZN(n368) );
  XNOR2_X1 U481 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n369) );
  XOR2_X1 U482 ( .A(n721), .B(n720), .Z(n370) );
  NOR2_X1 U483 ( .A1(n582), .A2(n372), .ZN(n605) );
  XNOR2_X1 U484 ( .A(n660), .B(KEYINPUT88), .ZN(n372) );
  XNOR2_X1 U485 ( .A(n465), .B(n464), .ZN(n724) );
  NOR2_X1 U486 ( .A1(n553), .A2(n693), .ZN(n513) );
  AND2_X2 U487 ( .A1(n543), .A2(n544), .ZN(n380) );
  NAND2_X1 U488 ( .A1(n512), .A2(n389), .ZN(n388) );
  INV_X1 U489 ( .A(n641), .ZN(n391) );
  NAND2_X1 U490 ( .A1(n625), .A2(n668), .ZN(n626) );
  INV_X1 U491 ( .A(n740), .ZN(n377) );
  NOR2_X1 U492 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U493 ( .A1(n550), .A2(n551), .ZN(n575) );
  NAND2_X1 U494 ( .A1(n378), .A2(n601), .ZN(n602) );
  NAND2_X1 U495 ( .A1(n593), .A2(n594), .ZN(n378) );
  AND2_X2 U496 ( .A1(n420), .A2(n617), .ZN(n751) );
  XNOR2_X2 U497 ( .A(n500), .B(n364), .ZN(n501) );
  OR2_X1 U498 ( .A1(n537), .A2(n368), .ZN(n409) );
  XNOR2_X1 U499 ( .A(n536), .B(KEYINPUT98), .ZN(n537) );
  XNOR2_X1 U500 ( .A(n381), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U501 ( .A1(n723), .A2(n737), .ZN(n381) );
  XNOR2_X1 U502 ( .A(n607), .B(n606), .ZN(n420) );
  NOR2_X2 U503 ( .A1(n692), .A2(n558), .ZN(n660) );
  NOR2_X2 U504 ( .A1(n570), .A2(n677), .ZN(n644) );
  XNOR2_X1 U505 ( .A(n447), .B(n382), .ZN(n448) );
  XNOR2_X2 U506 ( .A(n387), .B(n383), .ZN(n749) );
  XNOR2_X2 U507 ( .A(G143), .B(G128), .ZN(n447) );
  XNOR2_X2 U508 ( .A(n689), .B(n440), .ZN(n553) );
  XNOR2_X2 U509 ( .A(n384), .B(G472), .ZN(n689) );
  XNOR2_X2 U510 ( .A(n386), .B(n511), .ZN(n399) );
  NAND2_X1 U511 ( .A1(n628), .A2(n510), .ZN(n386) );
  XNOR2_X1 U512 ( .A(n387), .B(n394), .ZN(n476) );
  NOR2_X1 U513 ( .A1(n390), .A2(n393), .ZN(n392) );
  XNOR2_X2 U514 ( .A(n396), .B(KEYINPUT45), .ZN(n618) );
  XNOR2_X2 U515 ( .A(n398), .B(n400), .ZN(n397) );
  NAND2_X2 U516 ( .A1(n524), .A2(n527), .ZN(n398) );
  XNOR2_X2 U517 ( .A(n749), .B(G146), .ZN(n509) );
  NOR2_X1 U518 ( .A1(n693), .A2(n399), .ZN(n563) );
  XNOR2_X2 U519 ( .A(n403), .B(G122), .ZN(n469) );
  NAND2_X1 U520 ( .A1(n486), .A2(n533), .ZN(n487) );
  XNOR2_X2 U521 ( .A(n405), .B(n404), .ZN(n533) );
  XNOR2_X2 U522 ( .A(n556), .B(n481), .ZN(n583) );
  NAND2_X2 U523 ( .A1(n564), .A2(n674), .ZN(n556) );
  NAND2_X1 U524 ( .A1(n409), .A2(n407), .ZN(n406) );
  NAND2_X1 U525 ( .A1(n537), .A2(n408), .ZN(n407) );
  XNOR2_X2 U526 ( .A(n415), .B(n414), .ZN(n686) );
  XNOR2_X2 U527 ( .A(n501), .B(KEYINPUT77), .ZN(n415) );
  INV_X1 U528 ( .A(n569), .ZN(n675) );
  XNOR2_X1 U529 ( .A(n419), .B(n418), .ZN(n666) );
  NOR2_X1 U530 ( .A1(n760), .A2(n762), .ZN(n581) );
  XNOR2_X1 U531 ( .A(n428), .B(KEYINPUT121), .ZN(n716) );
  NAND2_X1 U532 ( .A1(n429), .A2(n431), .ZN(n428) );
  NAND2_X1 U533 ( .A1(n669), .A2(n668), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n722), .B(n370), .ZN(n723) );
  BUF_X1 U535 ( .A(n683), .Z(n712) );
  XNOR2_X2 U536 ( .A(n626), .B(KEYINPUT65), .ZN(n732) );
  XOR2_X1 U537 ( .A(n715), .B(KEYINPUT120), .Z(n431) );
  INV_X1 U538 ( .A(KEYINPUT68), .ZN(n522) );
  XNOR2_X1 U539 ( .A(n579), .B(KEYINPUT46), .ZN(n580) );
  XNOR2_X1 U540 ( .A(KEYINPUT48), .B(KEYINPUT87), .ZN(n606) );
  XNOR2_X1 U541 ( .A(n496), .B(n495), .ZN(n498) );
  INV_X1 U542 ( .A(n737), .ZN(n638) );
  XNOR2_X1 U543 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U544 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U545 ( .A1(G953), .A2(G237), .ZN(n455) );
  AND2_X1 U546 ( .A1(n455), .A2(G210), .ZN(n432) );
  XNOR2_X1 U547 ( .A(n432), .B(n471), .ZN(n438) );
  XNOR2_X1 U548 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U549 ( .A(KEYINPUT75), .B(KEYINPUT97), .ZN(n435) );
  XNOR2_X1 U550 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U551 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U552 ( .A(n509), .B(n439), .ZN(n634) );
  XNOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n440) );
  XOR2_X1 U554 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n444) );
  XNOR2_X2 U555 ( .A(n441), .B(KEYINPUT15), .ZN(n622) );
  INV_X1 U556 ( .A(n622), .ZN(n620) );
  NAND2_X1 U557 ( .A1(n620), .A2(G234), .ZN(n442) );
  XNOR2_X1 U558 ( .A(n442), .B(KEYINPUT20), .ZN(n499) );
  NAND2_X1 U559 ( .A1(G221), .A2(n499), .ZN(n443) );
  XNOR2_X1 U560 ( .A(n444), .B(n443), .ZN(n687) );
  XOR2_X1 U561 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n446) );
  XNOR2_X1 U562 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U563 ( .A(n448), .B(n470), .ZN(n449) );
  XOR2_X1 U564 ( .A(n450), .B(n449), .Z(n452) );
  NAND2_X1 U565 ( .A1(G217), .A2(n488), .ZN(n451) );
  XNOR2_X1 U566 ( .A(n452), .B(n451), .ZN(n729) );
  NOR2_X1 U567 ( .A1(G902), .A2(n729), .ZN(n453) );
  XNOR2_X1 U568 ( .A(G478), .B(n453), .ZN(n517) );
  AND2_X1 U569 ( .A1(n687), .A2(n517), .ZN(n467) );
  NAND2_X1 U570 ( .A1(G214), .A2(n455), .ZN(n456) );
  INV_X1 U571 ( .A(n457), .ZN(n458) );
  XOR2_X1 U572 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n462) );
  XNOR2_X1 U573 ( .A(G140), .B(KEYINPUT11), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n469), .B(KEYINPUT12), .ZN(n463) );
  NOR2_X1 U575 ( .A1(G902), .A2(n724), .ZN(n466) );
  NAND2_X1 U576 ( .A1(n467), .A2(n570), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n468), .B(KEYINPUT105), .ZN(n486) );
  XNOR2_X1 U578 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n481) );
  NAND2_X1 U579 ( .A1(G224), .A2(n752), .ZN(n472) );
  XNOR2_X1 U580 ( .A(KEYINPUT92), .B(KEYINPUT79), .ZN(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U582 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n739), .B(n477), .ZN(n719) );
  NOR2_X2 U584 ( .A1(n719), .A2(n622), .ZN(n479) );
  NAND2_X1 U585 ( .A1(G210), .A2(n480), .ZN(n478) );
  XNOR2_X2 U586 ( .A(n479), .B(n478), .ZN(n564) );
  NAND2_X1 U587 ( .A1(G214), .A2(n480), .ZN(n674) );
  NOR2_X1 U588 ( .A1(G898), .A2(n752), .ZN(n738) );
  NAND2_X1 U589 ( .A1(n738), .A2(G902), .ZN(n482) );
  NAND2_X1 U590 ( .A1(G952), .A2(n752), .ZN(n546) );
  NAND2_X1 U591 ( .A1(n482), .A2(n546), .ZN(n484) );
  NAND2_X1 U592 ( .A1(G234), .A2(G237), .ZN(n483) );
  XNOR2_X1 U593 ( .A(n483), .B(KEYINPUT14), .ZN(n670) );
  AND2_X1 U594 ( .A1(n484), .A2(n670), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n487), .B(KEYINPUT22), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G221), .A2(n488), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n497), .B(n505), .ZN(n750) );
  NAND2_X1 U600 ( .A1(n499), .A2(G217), .ZN(n500) );
  XNOR2_X1 U601 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U602 ( .A(n505), .B(n504), .Z(n507) );
  NAND2_X1 U603 ( .A1(G227), .A2(n752), .ZN(n506) );
  XNOR2_X1 U604 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U605 ( .A(n509), .B(n508), .ZN(n628) );
  INV_X1 U606 ( .A(G469), .ZN(n511) );
  INV_X1 U607 ( .A(n689), .ZN(n574) );
  NAND2_X1 U608 ( .A1(n513), .A2(n611), .ZN(n514) );
  XNOR2_X1 U609 ( .A(n514), .B(KEYINPUT33), .ZN(n683) );
  NAND2_X1 U610 ( .A1(n683), .A2(n533), .ZN(n516) );
  XNOR2_X1 U611 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n515) );
  XNOR2_X1 U612 ( .A(n516), .B(n515), .ZN(n519) );
  INV_X1 U613 ( .A(n570), .ZN(n678) );
  INV_X1 U614 ( .A(n517), .ZN(n677) );
  NAND2_X1 U615 ( .A1(n678), .A2(n677), .ZN(n595) );
  INV_X1 U616 ( .A(n595), .ZN(n518) );
  NAND2_X1 U617 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U618 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n521), .B(n520), .ZN(n525) );
  OR2_X2 U620 ( .A1(n525), .A2(KEYINPUT44), .ZN(n523) );
  XNOR2_X2 U621 ( .A(n523), .B(n522), .ZN(n524) );
  INV_X1 U622 ( .A(KEYINPUT89), .ZN(n526) );
  NAND2_X1 U623 ( .A1(n642), .A2(n526), .ZN(n528) );
  NAND2_X1 U624 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U625 ( .A1(n529), .A2(KEYINPUT44), .ZN(n544) );
  INV_X1 U626 ( .A(n693), .ZN(n530) );
  NAND2_X1 U627 ( .A1(n530), .A2(n393), .ZN(n531) );
  NOR2_X2 U628 ( .A1(n531), .A2(n692), .ZN(n699) );
  NAND2_X1 U629 ( .A1(n533), .A2(n699), .ZN(n532) );
  XNOR2_X2 U630 ( .A(n532), .B(KEYINPUT31), .ZN(n657) );
  INV_X1 U631 ( .A(n533), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n574), .A2(n563), .ZN(n534) );
  NOR2_X1 U633 ( .A1(n535), .A2(n534), .ZN(n646) );
  NOR2_X1 U634 ( .A1(n657), .A2(n646), .ZN(n536) );
  INV_X1 U635 ( .A(n644), .ZN(n566) );
  AND2_X1 U636 ( .A1(n570), .A2(n677), .ZN(n656) );
  INV_X1 U637 ( .A(n656), .ZN(n608) );
  NAND2_X1 U638 ( .A1(n566), .A2(n608), .ZN(n591) );
  INV_X1 U639 ( .A(n591), .ZN(n672) );
  NAND2_X1 U640 ( .A1(n379), .A2(n553), .ZN(n538) );
  OR2_X1 U641 ( .A1(n538), .A2(n611), .ZN(n539) );
  NOR2_X1 U642 ( .A1(n540), .A2(n539), .ZN(n643) );
  NAND2_X1 U643 ( .A1(n642), .A2(KEYINPUT44), .ZN(n541) );
  NAND2_X1 U644 ( .A1(n541), .A2(KEYINPUT89), .ZN(n542) );
  INV_X1 U645 ( .A(n687), .ZN(n549) );
  NOR2_X1 U646 ( .A1(G900), .A2(n752), .ZN(n545) );
  NAND2_X1 U647 ( .A1(n545), .A2(G902), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U649 ( .A1(n548), .A2(n670), .ZN(n561) );
  NOR2_X1 U650 ( .A1(n549), .A2(n561), .ZN(n551) );
  INV_X1 U651 ( .A(n686), .ZN(n550) );
  INV_X1 U652 ( .A(n575), .ZN(n552) );
  INV_X1 U653 ( .A(n553), .ZN(n554) );
  NAND2_X1 U654 ( .A1(n555), .A2(n554), .ZN(n610) );
  XNOR2_X1 U655 ( .A(n610), .B(KEYINPUT110), .ZN(n557) );
  NAND2_X1 U656 ( .A1(n689), .A2(n674), .ZN(n559) );
  XNOR2_X1 U657 ( .A(n559), .B(KEYINPUT30), .ZN(n560) );
  NOR2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n596) );
  INV_X1 U660 ( .A(n564), .ZN(n614) );
  NOR2_X1 U661 ( .A1(n596), .A2(n569), .ZN(n565) );
  XNOR2_X1 U662 ( .A(KEYINPUT39), .B(n565), .ZN(n609) );
  NOR2_X1 U663 ( .A1(n609), .A2(n566), .ZN(n568) );
  XNOR2_X1 U664 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n567) );
  XNOR2_X1 U665 ( .A(n568), .B(n567), .ZN(n760) );
  XNOR2_X1 U666 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n571) );
  XNOR2_X1 U667 ( .A(n571), .B(KEYINPUT41), .ZN(n572) );
  XNOR2_X1 U668 ( .A(n573), .B(n572), .ZN(n703) );
  INV_X1 U669 ( .A(KEYINPUT28), .ZN(n577) );
  XNOR2_X1 U670 ( .A(n577), .B(n576), .ZN(n578) );
  INV_X1 U671 ( .A(KEYINPUT64), .ZN(n579) );
  XNOR2_X1 U672 ( .A(n581), .B(n580), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U674 ( .A(KEYINPUT82), .B(n585), .ZN(n587) );
  NAND2_X1 U675 ( .A1(KEYINPUT47), .A2(n587), .ZN(n586) );
  XNOR2_X1 U676 ( .A(n586), .B(KEYINPUT84), .ZN(n589) );
  INV_X1 U677 ( .A(n587), .ZN(n653) );
  OR2_X1 U678 ( .A1(KEYINPUT74), .A2(n653), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n603) );
  OR2_X1 U680 ( .A1(KEYINPUT69), .A2(n672), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n590), .B(KEYINPUT47), .ZN(n594) );
  NAND2_X1 U682 ( .A1(KEYINPUT74), .A2(n653), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U685 ( .A1(n614), .A2(n597), .ZN(n652) );
  XOR2_X1 U686 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n598) );
  NOR2_X1 U687 ( .A1(n672), .A2(n598), .ZN(n599) );
  NOR2_X1 U688 ( .A1(KEYINPUT74), .A2(n599), .ZN(n600) );
  NOR2_X1 U689 ( .A1(n652), .A2(n600), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n607) );
  NOR2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n662) );
  NOR2_X1 U693 ( .A1(n390), .A2(n610), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n612), .A2(n674), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n663) );
  INV_X1 U697 ( .A(n663), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n662), .A2(n616), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n751), .ZN(n619) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n664) );
  NOR2_X1 U701 ( .A1(n620), .A2(KEYINPUT67), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(KEYINPUT2), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(KEYINPUT67), .ZN(n624) );
  INV_X1 U704 ( .A(n618), .ZN(n740) );
  NAND2_X1 U705 ( .A1(n732), .A2(G469), .ZN(n630) );
  XNOR2_X1 U706 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U709 ( .A1(n631), .A2(n737), .ZN(n633) );
  INV_X1 U710 ( .A(KEYINPUT123), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n633), .B(n632), .ZN(G54) );
  NAND2_X1 U712 ( .A1(n732), .A2(G472), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n634), .B(KEYINPUT62), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n636), .B(n635), .ZN(n637) );
  INV_X1 U715 ( .A(n637), .ZN(n639) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U718 ( .A(G110), .B(n641), .Z(G12) );
  XOR2_X1 U719 ( .A(n642), .B(G122), .Z(G24) );
  XOR2_X1 U720 ( .A(G101), .B(n643), .Z(G3) );
  NAND2_X1 U721 ( .A1(n646), .A2(n644), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n645), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n648) );
  NAND2_X1 U724 ( .A1(n646), .A2(n656), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U726 ( .A(G107), .B(n649), .ZN(G9) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U728 ( .A1(n656), .A2(n653), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(G30) );
  XOR2_X1 U730 ( .A(G143), .B(n652), .Z(G45) );
  NAND2_X1 U731 ( .A1(n653), .A2(n644), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(G146), .ZN(G48) );
  NAND2_X1 U733 ( .A1(n657), .A2(n644), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(G113), .ZN(G15) );
  XOR2_X1 U735 ( .A(G116), .B(KEYINPUT111), .Z(n659) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(G18) );
  XNOR2_X1 U738 ( .A(G125), .B(n660), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U740 ( .A(G134), .B(n662), .Z(G36) );
  XNOR2_X1 U741 ( .A(G140), .B(n663), .ZN(G42) );
  XOR2_X1 U742 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n718) );
  NAND2_X1 U743 ( .A1(n358), .A2(n664), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n667), .B(KEYINPUT83), .ZN(n669) );
  INV_X1 U746 ( .A(n670), .ZN(n710) );
  XNOR2_X1 U747 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n708) );
  NOR2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n673), .B(KEYINPUT117), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U751 ( .A(KEYINPUT116), .B(n676), .Z(n680) );
  NOR2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n684), .A2(n712), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT118), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n687), .A2(n379), .ZN(n688) );
  XOR2_X1 U758 ( .A(KEYINPUT49), .B(n688), .Z(n690) );
  NOR2_X1 U759 ( .A1(n690), .A2(n393), .ZN(n691) );
  XOR2_X1 U760 ( .A(n691), .B(KEYINPUT112), .Z(n697) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(KEYINPUT113), .ZN(n695) );
  XNOR2_X1 U763 ( .A(KEYINPUT50), .B(n695), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(KEYINPUT114), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U767 ( .A(n701), .B(KEYINPUT51), .Z(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT115), .B(n702), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U773 ( .A1(G952), .A2(n711), .ZN(n714) );
  NAND2_X1 U774 ( .A1(n703), .A2(n712), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U776 ( .A1(n716), .A2(n752), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n718), .B(n717), .ZN(G75) );
  NAND2_X1 U778 ( .A1(n732), .A2(G210), .ZN(n722) );
  XNOR2_X1 U779 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n721) );
  XNOR2_X1 U780 ( .A(n719), .B(KEYINPUT90), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n732), .A2(G475), .ZN(n726) );
  XOR2_X1 U782 ( .A(n724), .B(KEYINPUT59), .Z(n725) );
  XNOR2_X1 U783 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X2 U784 ( .A1(n727), .A2(n737), .ZN(n728) );
  XNOR2_X1 U785 ( .A(n728), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U786 ( .A1(n732), .A2(G478), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n729), .B(n730), .ZN(n731) );
  NOR2_X1 U788 ( .A1(n737), .A2(n731), .ZN(G63) );
  NAND2_X1 U789 ( .A1(n732), .A2(G217), .ZN(n735) );
  NOR2_X1 U790 ( .A1(n737), .A2(n736), .ZN(G66) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n748) );
  NOR2_X1 U792 ( .A1(n740), .A2(G953), .ZN(n741) );
  XOR2_X1 U793 ( .A(KEYINPUT126), .B(n741), .Z(n746) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U796 ( .A1(n743), .A2(G898), .ZN(n744) );
  XOR2_X1 U797 ( .A(KEYINPUT125), .B(n744), .Z(n745) );
  NAND2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n748), .B(n747), .ZN(G69) );
  XNOR2_X1 U800 ( .A(n749), .B(n750), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n751), .B(n754), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(n752), .ZN(n759) );
  XNOR2_X1 U803 ( .A(n754), .B(G227), .ZN(n755) );
  XNOR2_X1 U804 ( .A(n755), .B(KEYINPUT127), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n759), .A2(n758), .ZN(G72) );
  XOR2_X1 U808 ( .A(n760), .B(G131), .Z(G33) );
  XNOR2_X1 U809 ( .A(n761), .B(G119), .ZN(G21) );
  XOR2_X1 U810 ( .A(G137), .B(n762), .Z(G39) );
endmodule

