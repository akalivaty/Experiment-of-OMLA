

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U325 ( .A(n548), .B(KEYINPUT28), .Z(n512) );
  XNOR2_X1 U326 ( .A(G134GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U327 ( .A(n293), .B(KEYINPUT0), .ZN(n399) );
  XNOR2_X1 U328 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n294) );
  XNOR2_X1 U329 ( .A(n294), .B(KEYINPUT2), .ZN(n412) );
  XNOR2_X1 U330 ( .A(n399), .B(n412), .ZN(n313) );
  XOR2_X1 U331 ( .A(KEYINPUT4), .B(G57GAT), .Z(n296) );
  XNOR2_X1 U332 ( .A(G127GAT), .B(G148GAT), .ZN(n295) );
  XNOR2_X1 U333 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U334 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n298) );
  XNOR2_X1 U335 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n297) );
  XNOR2_X1 U336 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U337 ( .A(n300), .B(n299), .Z(n311) );
  XOR2_X1 U338 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n302) );
  XNOR2_X1 U339 ( .A(KEYINPUT6), .B(KEYINPUT87), .ZN(n301) );
  XNOR2_X1 U340 ( .A(n302), .B(n301), .ZN(n309) );
  XOR2_X1 U341 ( .A(G113GAT), .B(G1GAT), .Z(n324) );
  XOR2_X1 U342 ( .A(G85GAT), .B(G155GAT), .Z(n304) );
  XNOR2_X1 U343 ( .A(G29GAT), .B(G162GAT), .ZN(n303) );
  XNOR2_X1 U344 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U345 ( .A(n324), .B(n305), .Z(n307) );
  NAND2_X1 U346 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U348 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U349 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U350 ( .A(n313), .B(n312), .ZN(n546) );
  INV_X1 U351 ( .A(n546), .ZN(n471) );
  XOR2_X1 U352 ( .A(G15GAT), .B(G141GAT), .Z(n315) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(G197GAT), .ZN(n314) );
  XNOR2_X1 U354 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U355 ( .A(G8GAT), .B(KEYINPUT68), .Z(n317) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(KEYINPUT30), .ZN(n316) );
  XNOR2_X1 U357 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U358 ( .A(n319), .B(n318), .ZN(n329) );
  XOR2_X1 U359 ( .A(G29GAT), .B(G43GAT), .Z(n321) );
  XNOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U361 ( .A(n321), .B(n320), .ZN(n359) );
  XOR2_X1 U362 ( .A(n359), .B(KEYINPUT29), .Z(n323) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U364 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U365 ( .A(n325), .B(n324), .Z(n327) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U367 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U368 ( .A(n329), .B(n328), .ZN(n569) );
  XOR2_X1 U369 ( .A(G64GAT), .B(G92GAT), .Z(n331) );
  XNOR2_X1 U370 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U371 ( .A(n331), .B(n330), .ZN(n392) );
  XOR2_X1 U372 ( .A(KEYINPUT33), .B(n392), .Z(n333) );
  XOR2_X1 U373 ( .A(KEYINPUT70), .B(G148GAT), .Z(n416) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(n416), .ZN(n332) );
  XNOR2_X1 U375 ( .A(n333), .B(n332), .ZN(n339) );
  XOR2_X1 U376 ( .A(G85GAT), .B(KEYINPUT71), .Z(n335) );
  XNOR2_X1 U377 ( .A(G99GAT), .B(G106GAT), .ZN(n334) );
  XNOR2_X1 U378 ( .A(n335), .B(n334), .ZN(n358) );
  XOR2_X1 U379 ( .A(n358), .B(KEYINPUT31), .Z(n337) );
  NAND2_X1 U380 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U381 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U382 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT13), .Z(n341) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U385 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U386 ( .A(KEYINPUT69), .B(n342), .Z(n367) );
  XOR2_X1 U387 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U388 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U389 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U390 ( .A(n367), .B(n345), .ZN(n346) );
  XNOR2_X1 U391 ( .A(n347), .B(n346), .ZN(n574) );
  NOR2_X1 U392 ( .A1(n569), .A2(n574), .ZN(n457) );
  XOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n349) );
  XNOR2_X1 U394 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n348) );
  XNOR2_X1 U395 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U396 ( .A(G36GAT), .B(G190GAT), .Z(n387) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n350) );
  XNOR2_X1 U398 ( .A(n350), .B(G162GAT), .ZN(n425) );
  XOR2_X1 U399 ( .A(n387), .B(n425), .Z(n352) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U402 ( .A(n354), .B(n353), .ZN(n363) );
  XOR2_X1 U403 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n356) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U406 ( .A(n357), .B(KEYINPUT76), .Z(n361) );
  XNOR2_X1 U407 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U408 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U409 ( .A(n363), .B(n362), .ZN(n498) );
  INV_X1 U410 ( .A(n498), .ZN(n563) );
  XOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT81), .Z(n365) );
  XNOR2_X1 U412 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n364) );
  XNOR2_X1 U413 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U414 ( .A(n367), .B(n366), .ZN(n379) );
  XOR2_X1 U415 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n369) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G127GAT), .Z(n395) );
  XOR2_X1 U417 ( .A(G22GAT), .B(G155GAT), .Z(n417) );
  XNOR2_X1 U418 ( .A(n395), .B(n417), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U420 ( .A(KEYINPUT77), .B(G211GAT), .Z(n371) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(G183GAT), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n383) );
  XOR2_X1 U423 ( .A(KEYINPUT79), .B(n383), .Z(n373) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U426 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U427 ( .A(G1GAT), .B(G64GAT), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U429 ( .A(n379), .B(n378), .ZN(n578) );
  INV_X1 U430 ( .A(n578), .ZN(n500) );
  NOR2_X1 U431 ( .A1(n563), .A2(n500), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n380), .B(KEYINPUT16), .ZN(n442) );
  XOR2_X1 U433 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n385) );
  XOR2_X1 U434 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n382) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n413) );
  XNOR2_X1 U437 ( .A(n413), .B(n383), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U439 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n391) );
  XNOR2_X1 U443 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n396) );
  XOR2_X1 U445 ( .A(n396), .B(n392), .Z(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n542) );
  XOR2_X1 U447 ( .A(KEYINPUT27), .B(n542), .Z(n436) );
  XOR2_X1 U448 ( .A(n396), .B(n395), .Z(n398) );
  XNOR2_X1 U449 ( .A(G43GAT), .B(G99GAT), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n398), .B(n397), .ZN(n403) );
  XOR2_X1 U451 ( .A(n399), .B(G176GAT), .Z(n401) );
  NAND2_X1 U452 ( .A1(G227GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U454 ( .A(n403), .B(n402), .Z(n411) );
  XOR2_X1 U455 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n405) );
  XNOR2_X1 U456 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U458 ( .A(KEYINPUT20), .B(G71GAT), .Z(n407) );
  XNOR2_X1 U459 ( .A(G113GAT), .B(G183GAT), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n552) );
  INV_X1 U463 ( .A(n552), .ZN(n513) );
  XNOR2_X1 U464 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U465 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n415) );
  XNOR2_X1 U466 ( .A(G204GAT), .B(G78GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U468 ( .A(G211GAT), .B(G106GAT), .Z(n419) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U471 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U473 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U474 ( .A(n424), .B(KEYINPUT86), .Z(n427) );
  XNOR2_X1 U475 ( .A(n425), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U477 ( .A(n429), .B(n428), .ZN(n548) );
  NOR2_X1 U478 ( .A1(n513), .A2(n548), .ZN(n430) );
  XNOR2_X1 U479 ( .A(n430), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U480 ( .A1(n436), .A2(n567), .ZN(n434) );
  INV_X1 U481 ( .A(n542), .ZN(n488) );
  NAND2_X1 U482 ( .A1(n488), .A2(n513), .ZN(n431) );
  NAND2_X1 U483 ( .A1(n548), .A2(n431), .ZN(n432) );
  XOR2_X1 U484 ( .A(KEYINPUT25), .B(n432), .Z(n433) );
  NAND2_X1 U485 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U486 ( .A1(n435), .A2(n471), .ZN(n440) );
  NAND2_X1 U487 ( .A1(n436), .A2(n546), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n437), .B(KEYINPUT94), .ZN(n510) );
  NOR2_X1 U489 ( .A1(n512), .A2(n510), .ZN(n438) );
  NAND2_X1 U490 ( .A1(n552), .A2(n438), .ZN(n439) );
  NAND2_X1 U491 ( .A1(n440), .A2(n439), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT95), .B(n441), .Z(n453) );
  NAND2_X1 U493 ( .A1(n442), .A2(n453), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT96), .B(n443), .Z(n470) );
  NAND2_X1 U495 ( .A1(n457), .A2(n470), .ZN(n451) );
  NOR2_X1 U496 ( .A1(n471), .A2(n451), .ZN(n445) );
  XNOR2_X1 U497 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(G1GAT), .B(n446), .ZN(G1324GAT) );
  NOR2_X1 U500 ( .A1(n542), .A2(n451), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT98), .B(n447), .Z(n448) );
  XNOR2_X1 U502 ( .A(G8GAT), .B(n448), .ZN(G1325GAT) );
  NOR2_X1 U503 ( .A1(n552), .A2(n451), .ZN(n450) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(G1326GAT) );
  INV_X1 U506 ( .A(n512), .ZN(n477) );
  NOR2_X1 U507 ( .A1(n477), .A2(n451), .ZN(n452) );
  XOR2_X1 U508 ( .A(G22GAT), .B(n452), .Z(G1327GAT) );
  XOR2_X1 U509 ( .A(KEYINPUT38), .B(KEYINPUT100), .Z(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT36), .B(n498), .ZN(n583) );
  NAND2_X1 U511 ( .A1(n500), .A2(n453), .ZN(n454) );
  NOR2_X1 U512 ( .A1(n583), .A2(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(n483) );
  NAND2_X1 U515 ( .A1(n457), .A2(n483), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n467) );
  NAND2_X1 U517 ( .A1(n467), .A2(n546), .ZN(n462) );
  XNOR2_X1 U518 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT39), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(G1328GAT) );
  NAND2_X1 U521 ( .A1(n467), .A2(n488), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT102), .ZN(n464) );
  XNOR2_X1 U523 ( .A(G36GAT), .B(n464), .ZN(G1329GAT) );
  NAND2_X1 U524 ( .A1(n513), .A2(n467), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT40), .ZN(n466) );
  XNOR2_X1 U526 ( .A(G43GAT), .B(n466), .ZN(G1330GAT) );
  NAND2_X1 U527 ( .A1(n467), .A2(n512), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U529 ( .A(n574), .B(KEYINPUT41), .ZN(n517) );
  INV_X1 U530 ( .A(n517), .ZN(n555) );
  NAND2_X1 U531 ( .A1(n555), .A2(n569), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n469), .B(KEYINPUT103), .ZN(n484) );
  NAND2_X1 U533 ( .A1(n484), .A2(n470), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n471), .A2(n478), .ZN(n473) );
  XNOR2_X1 U535 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U537 ( .A(G57GAT), .B(n474), .Z(G1332GAT) );
  NOR2_X1 U538 ( .A1(n542), .A2(n478), .ZN(n475) );
  XOR2_X1 U539 ( .A(G64GAT), .B(n475), .Z(G1333GAT) );
  NOR2_X1 U540 ( .A1(n552), .A2(n478), .ZN(n476) );
  XOR2_X1 U541 ( .A(G71GAT), .B(n476), .Z(G1334GAT) );
  NOR2_X1 U542 ( .A1(n478), .A2(n477), .ZN(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n480) );
  XNOR2_X1 U544 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U545 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(G1335GAT) );
  NAND2_X1 U547 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(KEYINPUT107), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n492), .A2(n546), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n486), .B(KEYINPUT108), .ZN(n487) );
  XNOR2_X1 U551 ( .A(G85GAT), .B(n487), .ZN(G1336GAT) );
  NAND2_X1 U552 ( .A1(n492), .A2(n488), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n489), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U554 ( .A(G99GAT), .B(KEYINPUT109), .Z(n491) );
  NAND2_X1 U555 ( .A1(n492), .A2(n513), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(G1338GAT) );
  NAND2_X1 U557 ( .A1(n492), .A2(n512), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n493), .B(KEYINPUT44), .ZN(n494) );
  XNOR2_X1 U559 ( .A(G106GAT), .B(n494), .ZN(G1339GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT64), .B(KEYINPUT111), .Z(n509) );
  XNOR2_X1 U561 ( .A(n578), .B(KEYINPUT110), .ZN(n560) );
  NOR2_X1 U562 ( .A1(n569), .A2(n517), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n495), .B(KEYINPUT46), .ZN(n496) );
  NOR2_X1 U564 ( .A1(n560), .A2(n496), .ZN(n497) );
  NAND2_X1 U565 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n499), .B(KEYINPUT47), .ZN(n506) );
  NOR2_X1 U567 ( .A1(n500), .A2(n583), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(KEYINPUT45), .ZN(n502) );
  XNOR2_X1 U569 ( .A(KEYINPUT66), .B(n502), .ZN(n503) );
  NAND2_X1 U570 ( .A1(n503), .A2(n569), .ZN(n504) );
  NOR2_X1 U571 ( .A1(n504), .A2(n574), .ZN(n505) );
  NOR2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(KEYINPUT48), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n543) );
  NOR2_X1 U575 ( .A1(n543), .A2(n510), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(n511), .Z(n530) );
  NOR2_X1 U577 ( .A1(n512), .A2(n530), .ZN(n514) );
  NAND2_X1 U578 ( .A1(n514), .A2(n513), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n569), .A2(n522), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1340GAT) );
  NOR2_X1 U582 ( .A1(n522), .A2(n517), .ZN(n521) );
  XOR2_X1 U583 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n519) );
  XNOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n524) );
  INV_X1 U588 ( .A(n522), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n526), .A2(n560), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U591 ( .A(G127GAT), .B(n525), .Z(G1342GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n528) );
  NAND2_X1 U593 ( .A1(n526), .A2(n563), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(G134GAT), .B(n529), .Z(G1343GAT) );
  XNOR2_X1 U596 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n533) );
  INV_X1 U597 ( .A(n567), .ZN(n531) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n538) );
  INV_X1 U599 ( .A(n569), .ZN(n553) );
  NAND2_X1 U600 ( .A1(n538), .A2(n553), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  NAND2_X1 U603 ( .A1(n538), .A2(n555), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(G148GAT), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U606 ( .A1(n538), .A2(n578), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n537), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n540) );
  NAND2_X1 U609 ( .A1(n538), .A2(n563), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(G162GAT), .B(n541), .ZN(G1347GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n550) );
  NOR2_X1 U613 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U614 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n545), .B(n544), .ZN(n547) );
  NOR2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n568), .A2(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n553), .A2(n564), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT57), .Z(n557) );
  NAND2_X1 U623 ( .A1(n564), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n564), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n562), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n582), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n582), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

