

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U320 ( .A(n371), .B(n370), .Z(n554) );
  XNOR2_X1 U321 ( .A(n474), .B(n473), .ZN(n499) );
  XOR2_X1 U322 ( .A(n322), .B(n321), .Z(n519) );
  XNOR2_X1 U323 ( .A(n408), .B(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U324 ( .A(n309), .B(KEYINPUT93), .ZN(n310) );
  XNOR2_X1 U325 ( .A(n410), .B(n409), .ZN(n566) );
  XNOR2_X1 U326 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n405) );
  XNOR2_X1 U327 ( .A(n311), .B(n310), .ZN(n313) );
  XNOR2_X1 U328 ( .A(n406), .B(n405), .ZN(n543) );
  AND2_X1 U329 ( .A1(n528), .A2(n448), .ZN(n562) );
  XNOR2_X1 U330 ( .A(n353), .B(n352), .ZN(n571) );
  INV_X1 U331 ( .A(G36GAT), .ZN(n475) );
  XNOR2_X1 U332 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n449) );
  XNOR2_X1 U333 ( .A(n475), .B(KEYINPUT106), .ZN(n476) );
  XNOR2_X1 U334 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(n477), .B(n476), .ZN(G1329GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n289) );
  XNOR2_X1 U337 ( .A(G113GAT), .B(KEYINPUT66), .ZN(n288) );
  XNOR2_X1 U338 ( .A(n289), .B(n288), .ZN(n307) );
  XOR2_X1 U339 ( .A(G176GAT), .B(G190GAT), .Z(n291) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G99GAT), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U342 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n293) );
  XNOR2_X1 U343 ( .A(G71GAT), .B(G15GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U345 ( .A(n295), .B(n294), .Z(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT0), .B(G134GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G127GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(KEYINPUT81), .B(n298), .Z(n428) );
  XOR2_X1 U350 ( .A(G169GAT), .B(KEYINPUT19), .Z(n300) );
  XNOR2_X1 U351 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U353 ( .A(n308), .B(G183GAT), .Z(n302) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n428), .B(n303), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n521) );
  INV_X1 U359 ( .A(n521), .ZN(n528) );
  XNOR2_X1 U360 ( .A(KEYINPUT91), .B(n308), .ZN(n311) );
  AND2_X1 U361 ( .A1(G226GAT), .A2(G233GAT), .ZN(n309) );
  XOR2_X1 U362 ( .A(G190GAT), .B(G36GAT), .Z(n361) );
  XOR2_X1 U363 ( .A(n361), .B(KEYINPUT92), .Z(n312) );
  XOR2_X1 U364 ( .A(n313), .B(n312), .Z(n316) );
  XOR2_X1 U365 ( .A(G204GAT), .B(G176GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(G92GAT), .B(G64GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n336) );
  XNOR2_X1 U368 ( .A(n316), .B(n336), .ZN(n322) );
  XNOR2_X1 U369 ( .A(G183GAT), .B(G8GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n317), .B(KEYINPUT76), .ZN(n378) );
  XOR2_X1 U371 ( .A(KEYINPUT21), .B(G197GAT), .Z(n319) );
  XNOR2_X1 U372 ( .A(G218GAT), .B(KEYINPUT86), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(G211GAT), .B(n320), .Z(n442) );
  XNOR2_X1 U375 ( .A(n378), .B(n442), .ZN(n321) );
  INV_X1 U376 ( .A(n519), .ZN(n453) );
  XOR2_X1 U377 ( .A(n453), .B(KEYINPUT123), .Z(n407) );
  XNOR2_X1 U378 ( .A(G57GAT), .B(G71GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n323), .B(KEYINPUT13), .ZN(n372) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n324), .B(G78GAT), .ZN(n441) );
  XNOR2_X1 U382 ( .A(n372), .B(n441), .ZN(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n326) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n328) );
  INV_X1 U386 ( .A(KEYINPUT32), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n332) );
  INV_X1 U389 ( .A(KEYINPUT31), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U391 ( .A(G85GAT), .B(G99GAT), .Z(n362) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(n362), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(n336), .B(n335), .Z(n574) );
  INV_X1 U395 ( .A(n574), .ZN(n451) );
  XNOR2_X1 U396 ( .A(KEYINPUT70), .B(KEYINPUT7), .ZN(n337) );
  XNOR2_X1 U397 ( .A(n337), .B(KEYINPUT8), .ZN(n338) );
  XOR2_X1 U398 ( .A(n338), .B(KEYINPUT69), .Z(n340) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(G43GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n367) );
  XOR2_X1 U401 ( .A(G197GAT), .B(G169GAT), .Z(n342) );
  XNOR2_X1 U402 ( .A(G141GAT), .B(G22GAT), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n367), .B(n343), .ZN(n353) );
  XOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n345) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U408 ( .A(G15GAT), .B(KEYINPUT71), .Z(n383) );
  XOR2_X1 U409 ( .A(n383), .B(G50GAT), .Z(n347) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n421) );
  XNOR2_X1 U411 ( .A(n421), .B(G36GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U413 ( .A(n349), .B(n348), .Z(n351) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  INV_X1 U416 ( .A(KEYINPUT45), .ZN(n392) );
  XOR2_X1 U417 ( .A(G106GAT), .B(KEYINPUT74), .Z(n355) );
  XNOR2_X1 U418 ( .A(KEYINPUT9), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n371) );
  XOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT65), .Z(n357) );
  XNOR2_X1 U421 ( .A(G218GAT), .B(KEYINPUT67), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U423 ( .A(n358), .B(KEYINPUT11), .Z(n360) );
  XOR2_X1 U424 ( .A(G162GAT), .B(G50GAT), .Z(n433) );
  XNOR2_X1 U425 ( .A(G134GAT), .B(n433), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n366) );
  XOR2_X1 U427 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U430 ( .A(n366), .B(n365), .Z(n369) );
  XNOR2_X1 U431 ( .A(n367), .B(KEYINPUT10), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(KEYINPUT36), .B(n554), .ZN(n580) );
  XOR2_X1 U434 ( .A(n372), .B(KEYINPUT79), .Z(n377) );
  XOR2_X1 U435 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n374) );
  XNOR2_X1 U436 ( .A(KEYINPUT80), .B(KEYINPUT77), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n375), .B(KEYINPUT12), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n390) );
  XOR2_X1 U440 ( .A(G155GAT), .B(G22GAT), .Z(n432) );
  XOR2_X1 U441 ( .A(n432), .B(n378), .Z(n380) );
  NAND2_X1 U442 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U444 ( .A(G64GAT), .B(KEYINPUT14), .Z(n382) );
  XNOR2_X1 U445 ( .A(G211GAT), .B(G78GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U447 ( .A(n384), .B(n383), .Z(n386) );
  XNOR2_X1 U448 ( .A(G127GAT), .B(G1GAT), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U450 ( .A(n388), .B(n387), .Z(n389) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n478) );
  INV_X1 U452 ( .A(n478), .ZN(n577) );
  AND2_X1 U453 ( .A1(n580), .A2(n577), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U455 ( .A1(n571), .A2(n393), .ZN(n394) );
  NAND2_X1 U456 ( .A1(n451), .A2(n394), .ZN(n404) );
  XNOR2_X1 U457 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n395), .B(KEYINPUT47), .ZN(n402) );
  XOR2_X1 U459 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n396) );
  XOR2_X1 U461 ( .A(n396), .B(n574), .Z(n558) );
  NAND2_X1 U462 ( .A1(n571), .A2(n558), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n400) );
  NOR2_X1 U464 ( .A1(n577), .A2(n554), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  NAND2_X1 U467 ( .A1(n404), .A2(n403), .ZN(n406) );
  AND2_X1 U468 ( .A1(n407), .A2(n543), .ZN(n410) );
  INV_X1 U469 ( .A(KEYINPUT124), .ZN(n408) );
  XOR2_X1 U470 ( .A(G148GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U471 ( .A(G29GAT), .B(G85GAT), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U473 ( .A(G57GAT), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U474 ( .A(G155GAT), .B(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U476 ( .A(n416), .B(n415), .Z(n427) );
  XOR2_X1 U477 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n418) );
  XNOR2_X1 U478 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n425) );
  XOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT87), .Z(n420) );
  XNOR2_X1 U481 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n443) );
  XOR2_X1 U483 ( .A(n443), .B(n421), .Z(n423) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U488 ( .A(n429), .B(n428), .Z(n516) );
  XOR2_X1 U489 ( .A(KEYINPUT88), .B(KEYINPUT85), .Z(n431) );
  XNOR2_X1 U490 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n437) );
  XOR2_X1 U492 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n435) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U495 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U498 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n467) );
  NAND2_X1 U501 ( .A1(n516), .A2(n467), .ZN(n446) );
  OR2_X1 U502 ( .A1(n566), .A2(n446), .ZN(n447) );
  XNOR2_X1 U503 ( .A(KEYINPUT55), .B(n447), .ZN(n448) );
  NAND2_X1 U504 ( .A1(n562), .A2(n554), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n474) );
  NAND2_X1 U506 ( .A1(n451), .A2(n571), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n452), .B(KEYINPUT73), .ZN(n483) );
  XOR2_X1 U508 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n457) );
  NAND2_X1 U509 ( .A1(n528), .A2(n453), .ZN(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT97), .B(n454), .Z(n455) );
  NAND2_X1 U511 ( .A1(n455), .A2(n467), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n462) );
  XOR2_X1 U513 ( .A(n519), .B(KEYINPUT27), .Z(n465) );
  XNOR2_X1 U514 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT26), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n528), .A2(n467), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n546) );
  INV_X1 U518 ( .A(n546), .ZN(n568) );
  NAND2_X1 U519 ( .A1(n465), .A2(n568), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n463), .A2(n516), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT99), .ZN(n469) );
  INV_X1 U523 ( .A(n516), .ZN(n567) );
  AND2_X1 U524 ( .A1(n567), .A2(n465), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT94), .B(n466), .ZN(n544) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT28), .ZN(n525) );
  NAND2_X1 U527 ( .A1(n544), .A2(n525), .ZN(n530) );
  NOR2_X1 U528 ( .A1(n530), .A2(n528), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n481) );
  NOR2_X1 U530 ( .A1(n481), .A2(n577), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT104), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n580), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT37), .ZN(n515) );
  NAND2_X1 U534 ( .A1(n483), .A2(n515), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n499), .A2(n519), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n554), .A2(n478), .ZN(n479) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(n482), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n483), .A2(n504), .ZN(n491) );
  NOR2_X1 U541 ( .A1(n516), .A2(n491), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(n484), .Z(n485) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n519), .A2(n491), .ZN(n486) );
  XOR2_X1 U545 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U546 ( .A1(n491), .A2(n521), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n488) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n525), .A2(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n516), .A2(n499), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(KEYINPUT39), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n499), .A2(n521), .ZN(n497) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  INV_X1 U561 ( .A(KEYINPUT108), .ZN(n501) );
  NOR2_X1 U562 ( .A1(n499), .A2(n525), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  INV_X1 U565 ( .A(n558), .ZN(n503) );
  NOR2_X1 U566 ( .A1(n571), .A2(n503), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n514), .A2(n504), .ZN(n510) );
  NOR2_X1 U568 ( .A1(n516), .A2(n510), .ZN(n505) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(KEYINPUT42), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n519), .A2(n510), .ZN(n507) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n521), .A2(n510), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U576 ( .A1(n525), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n516), .A2(n524), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n524), .ZN(n520) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n524), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U593 ( .A1(n528), .A2(n543), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n539), .A2(n571), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U598 ( .A1(n539), .A2(n558), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n538) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n536) );
  NAND2_X1 U602 ( .A1(n539), .A2(n577), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n554), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT121), .Z(n548) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n555), .A2(n571), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n555), .A2(n558), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n577), .A2(n555), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n562), .A2(n571), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n577), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT60), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT59), .B(n565), .Z(n573) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT125), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

