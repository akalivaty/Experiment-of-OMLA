//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT79), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT79), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G155gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n204), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT81), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212));
  INV_X1    g011(.A(new_n208), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT79), .B(G155gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n212), .B(KEYINPUT2), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n211), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G155gat), .B(G162gat), .ZN(new_n222));
  XOR2_X1   g021(.A(G141gat), .B(G148gat), .Z(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n210), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n202), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G228gat), .A2(G233gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT75), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT22), .ZN(new_n234));
  OAI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(new_n231), .B2(new_n232), .ZN(new_n235));
  INV_X1    g034(.A(G204gat), .ZN(new_n236));
  INV_X1    g035(.A(G197gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n237), .A2(KEYINPUT74), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(KEYINPUT74), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT74), .B(G197gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G204gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT75), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n245), .A3(new_n240), .A4(new_n242), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n204), .A2(new_n206), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT80), .B(G162gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n210), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n220), .B1(new_n253), .B2(new_n212), .ZN(new_n254));
  INV_X1    g053(.A(new_n217), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n202), .B(new_n225), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n249), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n223), .A2(new_n222), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(KEYINPUT81), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n224), .B1(new_n260), .B2(new_n217), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(new_n250), .A3(new_n248), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n230), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(KEYINPUT86), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n247), .A2(new_n267), .A3(new_n250), .A4(new_n248), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n202), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n225), .B1(new_n254), .B2(new_n255), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n265), .B1(new_n271), .B2(new_n229), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(new_n262), .B2(KEYINPUT86), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n261), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  OAI211_X1 g073(.A(KEYINPUT87), .B(new_n228), .C1(new_n274), .C2(new_n257), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n264), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G22gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT88), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT31), .B(G50gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n276), .A2(new_n277), .ZN(new_n283));
  AOI211_X1 g082(.A(G22gat), .B(new_n264), .C1(new_n272), .C2(new_n275), .ZN(new_n284));
  OAI22_X1  g083(.A1(new_n278), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n272), .A2(new_n275), .ZN(new_n286));
  INV_X1    g085(.A(new_n264), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G22gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n276), .A2(new_n277), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(KEYINPUT88), .A3(new_n290), .A4(new_n281), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT0), .ZN(new_n294));
  XNOR2_X1  g093(.A(G57gat), .B(G85gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G134gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G127gat), .ZN(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G134gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G113gat), .A2(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT70), .B1(new_n303), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NOR2_X1   g109(.A1(G113gat), .A2(G120gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT69), .B1(new_n310), .B2(new_n311), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n306), .A2(new_n317), .A3(new_n307), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(new_n302), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n301), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT68), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n313), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n309), .B(new_n315), .C1(new_n320), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT82), .B1(new_n270), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n315), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n322), .A2(new_n324), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n261), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n270), .A2(KEYINPUT83), .A3(new_n326), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT83), .B1(new_n270), .B2(new_n326), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n327), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n335), .B2(new_n338), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n327), .A2(new_n332), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n261), .A2(new_n330), .A3(KEYINPUT4), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n256), .A2(new_n326), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n337), .C1(new_n344), .C2(new_n226), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT5), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n339), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n227), .A2(new_n326), .A3(new_n256), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n348), .A2(new_n337), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n327), .A2(new_n332), .A3(KEYINPUT4), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n261), .A2(new_n330), .A3(new_n352), .A4(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n329), .A2(new_n319), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n309), .A2(new_n315), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n221), .A2(new_n354), .A3(new_n225), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT85), .B1(new_n356), .B2(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n349), .A2(new_n350), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n297), .B1(new_n347), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n333), .A2(new_n334), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n327), .A2(new_n332), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n338), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT84), .ZN(new_n366));
  INV_X1    g165(.A(new_n345), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n327), .A2(new_n332), .A3(new_n341), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n350), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n296), .A3(new_n359), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(new_n362), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(KEYINPUT6), .B(new_n297), .C1(new_n347), .C2(new_n360), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  AND2_X1   g175(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT64), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT64), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G169gat), .ZN(new_n387));
  INV_X1    g186(.A(G176gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT23), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT25), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT66), .ZN(new_n395));
  OR2_X1    g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n397), .C1(new_n383), .C2(KEYINPUT65), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n381), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT25), .A4(new_n392), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n395), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n383), .A2(KEYINPUT65), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AND4_X1   g205(.A1(KEYINPUT25), .A2(new_n389), .A3(new_n391), .A4(new_n392), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT66), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n394), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT27), .B(G183gat), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n412), .A2(KEYINPUT28), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT67), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n387), .A3(new_n388), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n416), .A2(KEYINPUT26), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(KEYINPUT26), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n392), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT76), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n386), .A2(new_n393), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT66), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT66), .B1(new_n406), .B2(new_n407), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n420), .ZN(new_n430));
  INV_X1    g229(.A(G226gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT29), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n420), .A3(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(new_n249), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n428), .B2(new_n420), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n430), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n433), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n438), .B(KEYINPUT77), .C1(new_n442), .C2(new_n437), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT77), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n431), .B(new_n432), .C1(new_n422), .C2(new_n430), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n444), .B(new_n249), .C1(new_n445), .C2(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G8gat), .B(G36gat), .Z(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT78), .ZN(new_n449));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n446), .A3(new_n451), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(KEYINPUT30), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n447), .A2(new_n456), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n330), .B1(new_n409), .B2(new_n421), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n428), .A2(new_n326), .A3(new_n420), .ZN(new_n460));
  INV_X1    g259(.A(G227gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n432), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G15gat), .B(G43gat), .Z(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT71), .ZN(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT33), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n463), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n467), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n463), .B2(KEYINPUT32), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n460), .ZN(new_n482));
  INV_X1    g281(.A(new_n462), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g283(.A(KEYINPUT34), .B(new_n462), .C1(new_n459), .C2(new_n460), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n479), .A2(new_n480), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n486), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n471), .A2(new_n472), .B1(new_n477), .B2(new_n475), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(KEYINPUT73), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n292), .A2(new_n375), .A3(new_n458), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT35), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n479), .A2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n489), .A2(new_n486), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n285), .B2(new_n291), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n373), .A2(new_n374), .B1(new_n455), .B2(new_n457), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT36), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(new_n502), .A3(new_n496), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n372), .A2(new_n362), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n296), .B1(new_n371), .B2(new_n359), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n374), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n458), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n285), .A2(new_n291), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n337), .B1(new_n358), .B2(new_n348), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT89), .B(KEYINPUT39), .Z(new_n513));
  AOI21_X1  g312(.A(new_n297), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n327), .A2(new_n332), .A3(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n357), .A2(new_n353), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n348), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n338), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  INV_X1    g318(.A(new_n335), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n337), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT40), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n506), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n514), .A2(new_n522), .A3(KEYINPUT40), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n524), .A2(new_n457), .A3(new_n455), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n447), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n435), .A2(new_n249), .A3(new_n436), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(KEYINPUT37), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n437), .B1(new_n445), .B2(new_n440), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n451), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n373), .A2(new_n374), .A3(new_n535), .A4(new_n453), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n452), .B1(new_n447), .B2(new_n527), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n443), .A2(new_n446), .A3(KEYINPUT37), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n292), .B(new_n526), .C1(new_n536), .C2(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n493), .A2(new_n500), .B1(new_n511), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G197gat), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT11), .B(G169gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT12), .Z(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(KEYINPUT94), .C1(G1gat), .C2(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  INV_X1    g353(.A(G43gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(G50gat), .ZN(new_n556));
  INV_X1    g355(.A(G50gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(G43gat), .B2(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n554), .A2(new_n555), .A3(G50gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT15), .B1(new_n555), .B2(G50gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n555), .B2(G50gat), .ZN(new_n562));
  INV_X1    g361(.A(G29gat), .ZN(new_n563));
  INV_X1    g362(.A(G36gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT14), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT91), .ZN(new_n573));
  INV_X1    g372(.A(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n560), .A2(new_n570), .B1(new_n575), .B2(new_n562), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n560), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n562), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT17), .B1(new_n582), .B2(KEYINPUT93), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n552), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n550), .B(G8gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n582), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT18), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(G229gat), .B2(G233gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n552), .A2(new_n576), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT13), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n552), .A2(new_n576), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n578), .B1(new_n576), .B2(new_n577), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n599), .B2(new_n552), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT18), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n546), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n592), .A3(new_n586), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n587), .ZN(new_n604));
  INV_X1    g403(.A(new_n546), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n604), .A2(new_n594), .A3(new_n589), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n606), .A3(KEYINPUT95), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n546), .C1(new_n595), .C2(new_n601), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT96), .B1(new_n607), .B2(new_n609), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G57gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G64gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT9), .ZN(new_n622));
  NAND2_X1  g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT97), .B1(G71gat), .B2(G78gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n623), .ZN(new_n626));
  NOR3_X1   g425(.A1(KEYINPUT97), .A2(G71gat), .A3(G78gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G57gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(G64gat), .ZN(new_n630));
  INV_X1    g429(.A(G64gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT9), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n620), .A2(new_n624), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n585), .B1(KEYINPUT21), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n203), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n634), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G127gat), .ZN(new_n643));
  XOR2_X1   g442(.A(G183gat), .B(G211gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  INV_X1    g446(.A(G85gat), .ZN(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT7), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT7), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n647), .B(new_n653), .C1(new_n648), .C2(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(G99gat), .A2(G106gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(KEYINPUT8), .A2(new_n655), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G99gat), .B(G106gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n660), .A2(new_n652), .A3(new_n654), .A4(new_n656), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT100), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n582), .A2(new_n662), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT102), .ZN(new_n667));
  INV_X1    g466(.A(new_n661), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n657), .A2(new_n658), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n599), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n667), .B2(new_n670), .ZN(new_n674));
  XNOR2_X1  g473(.A(G190gat), .B(G218gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G134gat), .B(G162gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n673), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n673), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n646), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n620), .A2(new_n624), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n628), .A2(new_n633), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n669), .B2(new_n668), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT10), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n659), .A2(new_n634), .A3(new_n661), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n689), .B2(new_n688), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n662), .A2(KEYINPUT103), .A3(KEYINPUT10), .A4(new_n634), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(G230gat), .A2(G233gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n687), .A2(new_n689), .ZN(new_n697));
  INV_X1    g496(.A(new_n695), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(G120gat), .B(G148gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(G176gat), .B(G204gat), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n701), .B(new_n702), .Z(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n683), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n541), .A2(new_n617), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n375), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  INV_X1    g512(.A(new_n458), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT16), .B(G8gat), .Z(new_n715));
  AND3_X1   g514(.A1(new_n710), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n551), .B1(new_n710), .B2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(KEYINPUT42), .B2(new_n716), .ZN(G1325gat));
  INV_X1    g518(.A(G15gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n494), .A2(new_n496), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n710), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n710), .A2(new_n504), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n720), .ZN(G1326gat));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n510), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  NOR2_X1   g527(.A1(new_n541), .A2(new_n617), .ZN(new_n729));
  INV_X1    g528(.A(new_n646), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n681), .A3(new_n707), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n563), .A3(new_n711), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n541), .B2(new_n681), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n501), .A2(new_n503), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n499), .B2(new_n292), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n536), .A2(new_n539), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n526), .A2(new_n292), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n492), .A2(KEYINPUT35), .B1(new_n499), .B2(new_n498), .ZN(new_n743));
  OAI211_X1 g542(.A(KEYINPUT44), .B(new_n682), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n610), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n745), .A2(new_n746), .A3(new_n646), .A4(new_n708), .ZN(new_n747));
  OAI21_X1  g546(.A(G29gat), .B1(new_n747), .B2(new_n375), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n735), .A2(new_n748), .ZN(G1328gat));
  OAI21_X1  g548(.A(G36gat), .B1(new_n747), .B2(new_n458), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n732), .A2(G36gat), .A3(new_n458), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(G1329gat));
  OAI21_X1  g557(.A(G43gat), .B1(new_n747), .B2(new_n738), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n733), .A2(new_n555), .A3(new_n722), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT47), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n759), .B(new_n760), .C1(new_n762), .C2(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1330gat));
  OAI21_X1  g565(.A(new_n557), .B1(new_n732), .B2(new_n292), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n510), .A2(G50gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n747), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n683), .A2(new_n610), .A3(new_n707), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n541), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n541), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n375), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n629), .ZN(G1332gat));
  INV_X1    g576(.A(new_n775), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n714), .B1(new_n779), .B2(new_n631), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n631), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  OAI21_X1  g583(.A(G71gat), .B1(new_n775), .B2(new_n738), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n721), .A2(G71gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n775), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n778), .A2(new_n510), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n541), .A2(new_n681), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n730), .A2(new_n746), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT51), .ZN(new_n795));
  NOR4_X1   g594(.A1(new_n795), .A2(G85gat), .A3(new_n375), .A4(new_n708), .ZN(new_n796));
  INV_X1    g595(.A(new_n793), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n708), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n745), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n648), .B1(new_n799), .B2(new_n711), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n796), .A2(new_n800), .ZN(G1336gat));
  NAND4_X1  g600(.A1(new_n737), .A2(new_n714), .A3(new_n744), .A4(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n493), .A2(new_n500), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n511), .A2(new_n540), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n682), .A4(new_n793), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n811), .B2(KEYINPUT111), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT110), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n792), .B2(new_n793), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n714), .A2(new_n649), .A3(new_n707), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n805), .B(new_n806), .C1(new_n816), .C2(KEYINPUT112), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n812), .A2(new_n814), .A3(new_n818), .A4(new_n815), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n803), .C1(new_n795), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1337gat));
  NOR4_X1   g622(.A1(new_n795), .A2(G99gat), .A3(new_n721), .A4(new_n708), .ZN(new_n824));
  INV_X1    g623(.A(G99gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n799), .B2(new_n504), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n824), .A2(new_n826), .ZN(G1338gat));
  NAND4_X1  g626(.A1(new_n737), .A2(new_n510), .A3(new_n744), .A4(new_n798), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G106gat), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n812), .A2(new_n814), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n292), .A2(G106gat), .A3(new_n708), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n829), .A2(new_n830), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n829), .B(new_n838), .C1(new_n795), .C2(new_n834), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1339gat));
  NAND3_X1  g639(.A1(new_n683), .A2(new_n610), .A3(new_n708), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n690), .A2(new_n693), .A3(new_n692), .A4(new_n698), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n696), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n694), .A2(new_n844), .A3(new_n695), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n843), .A2(KEYINPUT55), .A3(new_n704), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n706), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n704), .A3(new_n845), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n591), .A2(new_n593), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n600), .A2(new_n592), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n545), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n606), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n682), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n607), .A2(new_n847), .A3(new_n609), .A4(new_n850), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n606), .A3(new_n707), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n682), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(KEYINPUT116), .A3(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n841), .B1(new_n865), .B2(new_n730), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n866), .B2(new_n292), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n861), .A2(new_n862), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n681), .A3(new_n864), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n730), .B1(new_n870), .B2(new_n857), .ZN(new_n871));
  INV_X1    g670(.A(new_n841), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT117), .B(new_n292), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n711), .A3(new_n458), .A4(new_n722), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n617), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n866), .A2(new_n711), .A3(new_n292), .A4(new_n491), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n714), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n304), .B(new_n746), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n881), .ZN(G1340gat));
  OAI21_X1  g681(.A(G120gat), .B1(new_n875), .B2(new_n708), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n305), .B(new_n707), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n875), .B2(new_n646), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n300), .A3(new_n730), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1342gat));
  OAI21_X1  g687(.A(G134gat), .B1(new_n875), .B2(new_n681), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n877), .A2(G134gat), .A3(new_n714), .A4(new_n681), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n510), .A2(new_n738), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT121), .Z(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n866), .A3(new_n711), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n714), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n617), .A2(G141gat), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT58), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n711), .A2(new_n738), .A3(new_n458), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT119), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n866), .B2(new_n510), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n510), .A2(KEYINPUT57), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n851), .B1(new_n612), .B2(new_n614), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n682), .B1(new_n904), .B2(new_n860), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n646), .B1(new_n905), .B2(new_n858), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n841), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n901), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n899), .B1(new_n908), .B2(new_n617), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n908), .A2(new_n899), .A3(new_n617), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n898), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT120), .B(new_n901), .C1(new_n902), .C2(new_n907), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n746), .A3(new_n915), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n916), .A2(G141gat), .B1(new_n896), .B2(new_n897), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G1344gat));
  INV_X1    g718(.A(G148gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n914), .A2(new_n915), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n708), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n901), .A2(new_n707), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n906), .B1(new_n616), .B2(new_n709), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n925), .B2(new_n510), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n866), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n903), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n924), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT59), .B1(new_n931), .B2(new_n920), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n896), .A2(new_n920), .A3(new_n707), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(new_n251), .B1(new_n922), .B2(new_n646), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n896), .A2(new_n216), .A3(new_n730), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(new_n252), .B1(new_n922), .B2(new_n681), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n458), .A2(new_n682), .A3(new_n215), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n895), .B2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n928), .A2(new_n711), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n292), .A2(new_n714), .A3(new_n491), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n746), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n711), .A2(new_n458), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n721), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n874), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n617), .A2(new_n387), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G1348gat));
  NAND3_X1  g751(.A1(new_n945), .A2(new_n388), .A3(new_n707), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n950), .A2(new_n707), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n388), .ZN(G1349gat));
  NAND3_X1  g754(.A1(new_n874), .A2(new_n730), .A3(new_n949), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G183gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n945), .A2(new_n410), .A3(new_n730), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n957), .A2(new_n959), .A3(new_n958), .A4(new_n962), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n945), .A2(new_n411), .A3(new_n682), .ZN(new_n967));
  INV_X1    g766(.A(new_n873), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n682), .B(new_n949), .C1(new_n968), .C2(new_n867), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(G190gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n969), .B2(G190gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(KEYINPUT125), .B(new_n967), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1351gat));
  NOR2_X1   g776(.A1(new_n893), .A2(new_n458), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n942), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n237), .A3(new_n746), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n948), .A2(new_n504), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n926), .B2(new_n929), .ZN(new_n984));
  OAI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n617), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n982), .A2(new_n985), .ZN(G1352gat));
  AOI21_X1  g785(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n980), .A2(new_n707), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n988), .B(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(G204gat), .B1(new_n984), .B2(new_n708), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n980), .A2(new_n231), .A3(new_n730), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n730), .B(new_n983), .C1(new_n926), .C2(new_n929), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n984), .B2(new_n681), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n232), .A3(new_n682), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


