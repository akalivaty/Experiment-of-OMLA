

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n794), .A2(n793), .ZN(n811) );
  AND2_X1 U553 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X2 U554 ( .A1(n543), .A2(n542), .ZN(G160) );
  BUF_X2 U555 ( .A(n887), .Z(n516) );
  XOR2_X1 U556 ( .A(KEYINPUT17), .B(n536), .Z(n887) );
  INV_X1 U557 ( .A(KEYINPUT101), .ZN(n746) );
  XNOR2_X1 U558 ( .A(n677), .B(KEYINPUT88), .ZN(n786) );
  NAND2_X1 U559 ( .A1(G160), .A2(G40), .ZN(n677) );
  OR2_X1 U560 ( .A1(n791), .A2(n790), .ZN(n517) );
  NOR2_X1 U561 ( .A1(n932), .A2(n705), .ZN(n707) );
  XNOR2_X1 U562 ( .A(n730), .B(KEYINPUT97), .ZN(n726) );
  NAND2_X1 U563 ( .A1(n678), .A2(n785), .ZN(n679) );
  NAND2_X1 U564 ( .A1(n792), .A2(n517), .ZN(n793) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NOR2_X1 U566 ( .A1(G651), .A2(n638), .ZN(n650) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U568 ( .A(G651), .ZN(n523) );
  NOR2_X1 U569 ( .A1(n638), .A2(n523), .ZN(n642) );
  NAND2_X1 U570 ( .A1(n642), .A2(G76), .ZN(n518) );
  XNOR2_X1 U571 ( .A(KEYINPUT80), .B(n518), .ZN(n521) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U573 ( .A1(n641), .A2(G89), .ZN(n519) );
  XNOR2_X1 U574 ( .A(KEYINPUT4), .B(n519), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U576 ( .A(KEYINPUT5), .B(n522), .ZN(n531) );
  NOR2_X1 U577 ( .A1(G543), .A2(n523), .ZN(n525) );
  XNOR2_X1 U578 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n524) );
  XNOR2_X1 U579 ( .A(n525), .B(n524), .ZN(n646) );
  NAND2_X1 U580 ( .A1(n646), .A2(G63), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT81), .B(n526), .Z(n528) );
  NAND2_X1 U582 ( .A1(n650), .A2(G51), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U584 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U586 ( .A(KEYINPUT7), .B(n532), .ZN(G168) );
  AND2_X1 U587 ( .A1(G2104), .A2(G101), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n534), .B(KEYINPUT65), .ZN(n535) );
  XNOR2_X1 U590 ( .A(n535), .B(KEYINPUT23), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G137), .A2(n516), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n543) );
  AND2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U594 ( .A1(G113), .A2(n883), .ZN(n541) );
  INV_X1 U595 ( .A(G2105), .ZN(n539) );
  NOR2_X2 U596 ( .A1(G2104), .A2(n539), .ZN(n881) );
  NAND2_X1 U597 ( .A1(G125), .A2(n881), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G64), .A2(n646), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G52), .A2(n650), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n642), .A2(G77), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT69), .B(n546), .Z(n548) );
  NAND2_X1 U604 ( .A1(n641), .A2(G90), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U607 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(G88), .A2(n641), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G75), .A2(n642), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G62), .A2(n646), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G50), .A2(n650), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(G166) );
  NAND2_X1 U618 ( .A1(n516), .A2(G138), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G114), .A2(n883), .ZN(n558) );
  XOR2_X1 U620 ( .A(KEYINPUT87), .B(n558), .Z(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G126), .A2(n881), .ZN(n562) );
  AND2_X1 U623 ( .A1(n539), .A2(G2104), .ZN(n888) );
  NAND2_X1 U624 ( .A1(G102), .A2(n888), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U626 ( .A1(n564), .A2(n563), .ZN(G164) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(n565) );
  XNOR2_X1 U628 ( .A(KEYINPUT82), .B(n565), .ZN(G286) );
  NAND2_X1 U629 ( .A1(G94), .A2(G452), .ZN(n566) );
  XOR2_X1 U630 ( .A(KEYINPUT70), .B(n566), .Z(G173) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n569) );
  INV_X1 U634 ( .A(G223), .ZN(n830) );
  NAND2_X1 U635 ( .A1(G567), .A2(n830), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G234) );
  XNOR2_X1 U637 ( .A(KEYINPUT75), .B(KEYINPUT13), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G81), .A2(n641), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT74), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G68), .A2(n642), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G56), .A2(n646), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT14), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT73), .ZN(n578) );
  NOR2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT76), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G43), .A2(n650), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n949) );
  INV_X1 U651 ( .A(G860), .ZN(n620) );
  OR2_X1 U652 ( .A1(n949), .A2(n620), .ZN(G153) );
  XNOR2_X1 U653 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G92), .A2(n641), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT78), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G66), .A2(n646), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G54), .A2(n650), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G79), .A2(n642), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT79), .B(n586), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U664 ( .A(KEYINPUT15), .B(n591), .ZN(n943) );
  OR2_X1 U665 ( .A1(n943), .A2(G868), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G65), .A2(n646), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G53), .A2(n650), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G91), .A2(n641), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G78), .A2(n642), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U675 ( .A1(G868), .A2(G286), .ZN(n602) );
  INV_X1 U676 ( .A(G299), .ZN(n932) );
  OR2_X1 U677 ( .A1(n932), .A2(G868), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n620), .A2(G559), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n603), .A2(n943), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n604), .B(KEYINPUT83), .ZN(n605) );
  XOR2_X1 U682 ( .A(KEYINPUT16), .B(n605), .Z(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n949), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G868), .A2(n943), .ZN(n606) );
  NOR2_X1 U685 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n881), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G135), .A2(n516), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G99), .A2(n888), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n883), .A2(G111), .ZN(n612) );
  XOR2_X1 U693 ( .A(KEYINPUT84), .B(n612), .Z(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n998) );
  XOR2_X1 U696 ( .A(n998), .B(G2096), .Z(n618) );
  XNOR2_X1 U697 ( .A(G2100), .B(KEYINPUT85), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n943), .ZN(n619) );
  XOR2_X1 U700 ( .A(n949), .B(n619), .Z(n658) );
  NAND2_X1 U701 ( .A1(n620), .A2(n658), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G67), .A2(n646), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G55), .A2(n650), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G93), .A2(n641), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G80), .A2(n642), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n661) );
  XOR2_X1 U709 ( .A(n627), .B(n661), .Z(G145) );
  NAND2_X1 U710 ( .A1(G86), .A2(n641), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G61), .A2(n646), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n642), .A2(G73), .ZN(n630) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n650), .A2(G48), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n650), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U721 ( .A1(n646), .A2(n637), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G85), .A2(n641), .ZN(n644) );
  NAND2_X1 U725 ( .A1(G72), .A2(n642), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U727 ( .A(KEYINPUT66), .B(n645), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n646), .A2(G60), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT68), .B(n647), .Z(n648) );
  NOR2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n650), .A2(G47), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(G290) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(G305), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(G288), .ZN(n654) );
  XOR2_X1 U735 ( .A(n654), .B(n661), .Z(n656) );
  XNOR2_X1 U736 ( .A(n932), .B(G166), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n657), .B(G290), .ZN(n900) );
  XNOR2_X1 U739 ( .A(n900), .B(n658), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n659), .A2(G868), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(KEYINPUT86), .ZN(n663) );
  OR2_X1 U742 ( .A1(G868), .A2(n661), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U752 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(G96), .A2(n670), .ZN(n834) );
  NAND2_X1 U754 ( .A1(n834), .A2(G2106), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G108), .A2(n672), .ZN(n835) );
  NAND2_X1 U758 ( .A1(n835), .A2(G567), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n836) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n836), .A2(n675), .ZN(n833) );
  NAND2_X1 U762 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U764 ( .A(G1981), .B(G305), .ZN(n951) );
  INV_X1 U765 ( .A(n786), .ZN(n678) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n785) );
  XNOR2_X1 U767 ( .A(n679), .B(KEYINPUT64), .ZN(n715) );
  BUF_X1 U768 ( .A(n715), .Z(n683) );
  NOR2_X1 U769 ( .A1(n683), .A2(G2084), .ZN(n716) );
  NAND2_X1 U770 ( .A1(n716), .A2(G8), .ZN(n728) );
  XNOR2_X1 U771 ( .A(G2078), .B(KEYINPUT92), .ZN(n680) );
  XNOR2_X1 U772 ( .A(n680), .B(KEYINPUT25), .ZN(n916) );
  INV_X1 U773 ( .A(n715), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n916), .A2(n700), .ZN(n682) );
  INV_X1 U775 ( .A(G1961), .ZN(n975) );
  NAND2_X1 U776 ( .A1(n683), .A2(n975), .ZN(n681) );
  NAND2_X1 U777 ( .A1(n682), .A2(n681), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n714), .A2(G171), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n683), .A2(G1341), .ZN(n687) );
  INV_X1 U780 ( .A(G1996), .ZN(n912) );
  NOR2_X1 U781 ( .A1(n715), .A2(n912), .ZN(n685) );
  XOR2_X1 U782 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n684) );
  XNOR2_X1 U783 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U784 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U785 ( .A1(n949), .A2(n688), .ZN(n691) );
  NOR2_X1 U786 ( .A1(n691), .A2(n943), .ZN(n690) );
  INV_X1 U787 ( .A(KEYINPUT96), .ZN(n689) );
  XNOR2_X1 U788 ( .A(n690), .B(n689), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n691), .A2(n943), .ZN(n696) );
  AND2_X1 U790 ( .A1(n700), .A2(G2067), .ZN(n692) );
  XNOR2_X1 U791 ( .A(n692), .B(KEYINPUT95), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n683), .A2(G1348), .ZN(n693) );
  NAND2_X1 U793 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G2072), .A2(n700), .ZN(n699) );
  XNOR2_X1 U797 ( .A(n699), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U798 ( .A(G1956), .ZN(n966) );
  NOR2_X1 U799 ( .A1(n700), .A2(n966), .ZN(n701) );
  NOR2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n932), .A2(n705), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n709) );
  XNOR2_X1 U803 ( .A(KEYINPUT28), .B(KEYINPUT93), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U806 ( .A(KEYINPUT29), .B(n710), .ZN(n711) );
  INV_X1 U807 ( .A(n711), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n724) );
  NOR2_X1 U809 ( .A1(G171), .A2(n714), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n715), .A2(G8), .ZN(n791) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n791), .ZN(n725) );
  NOR2_X1 U812 ( .A1(n725), .A2(n716), .ZN(n717) );
  NAND2_X1 U813 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U814 ( .A(n718), .B(KEYINPUT30), .ZN(n719) );
  NOR2_X1 U815 ( .A1(n719), .A2(G168), .ZN(n720) );
  NOR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(n722), .Z(n723) );
  NAND2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n743) );
  XNOR2_X1 U821 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n741) );
  AND2_X1 U822 ( .A1(G286), .A2(G8), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n739) );
  INV_X1 U824 ( .A(G8), .ZN(n737) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n791), .ZN(n731) );
  XNOR2_X1 U826 ( .A(n731), .B(KEYINPUT98), .ZN(n733) );
  NOR2_X1 U827 ( .A1(n683), .A2(G2090), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n734), .A2(G303), .ZN(n735) );
  XOR2_X1 U830 ( .A(KEYINPUT99), .B(n735), .Z(n736) );
  OR2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n760) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n937) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n937), .A2(n744), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n760), .A2(n745), .ZN(n747) );
  XNOR2_X1 U838 ( .A(n747), .B(n746), .ZN(n751) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n938) );
  INV_X1 U840 ( .A(n938), .ZN(n748) );
  NOR2_X1 U841 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  INV_X1 U842 ( .A(n791), .ZN(n752) );
  AND2_X1 U843 ( .A1(n749), .A2(n752), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n937), .A2(n752), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U848 ( .A(KEYINPUT102), .B(n756), .Z(n757) );
  NOR2_X1 U849 ( .A1(n951), .A2(n757), .ZN(n794) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U851 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n791), .A2(n761), .ZN(n788) );
  NAND2_X1 U854 ( .A1(G105), .A2(n888), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n762), .B(KEYINPUT38), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G141), .A2(n516), .ZN(n763) );
  XOR2_X1 U857 ( .A(KEYINPUT91), .B(n763), .Z(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U859 ( .A1(G117), .A2(n883), .ZN(n767) );
  NAND2_X1 U860 ( .A1(G129), .A2(n881), .ZN(n766) );
  NAND2_X1 U861 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U862 ( .A1(n769), .A2(n768), .ZN(n862) );
  AND2_X1 U863 ( .A1(n912), .A2(n862), .ZN(n993) );
  XOR2_X1 U864 ( .A(KEYINPUT90), .B(G1991), .Z(n917) );
  NAND2_X1 U865 ( .A1(n516), .A2(G131), .ZN(n772) );
  NAND2_X1 U866 ( .A1(G107), .A2(n883), .ZN(n770) );
  XOR2_X1 U867 ( .A(KEYINPUT89), .B(n770), .Z(n771) );
  NAND2_X1 U868 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U869 ( .A1(G119), .A2(n881), .ZN(n774) );
  NAND2_X1 U870 ( .A1(G95), .A2(n888), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n872) );
  AND2_X1 U873 ( .A1(n917), .A2(n872), .ZN(n1001) );
  NOR2_X1 U874 ( .A1(G1986), .A2(G290), .ZN(n777) );
  XOR2_X1 U875 ( .A(n777), .B(KEYINPUT103), .Z(n778) );
  NOR2_X1 U876 ( .A1(n1001), .A2(n778), .ZN(n782) );
  NOR2_X1 U877 ( .A1(n917), .A2(n872), .ZN(n780) );
  NOR2_X1 U878 ( .A1(n862), .A2(n912), .ZN(n779) );
  NOR2_X1 U879 ( .A1(n780), .A2(n779), .ZN(n1004) );
  INV_X1 U880 ( .A(n1004), .ZN(n781) );
  NOR2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U882 ( .A1(n993), .A2(n783), .ZN(n784) );
  XNOR2_X1 U883 ( .A(KEYINPUT39), .B(n784), .ZN(n787) );
  NOR2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n814) );
  NAND2_X1 U885 ( .A1(n787), .A2(n814), .ZN(n804) );
  AND2_X1 U886 ( .A1(n788), .A2(n804), .ZN(n792) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U888 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  XNOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NAND2_X1 U890 ( .A1(G140), .A2(n516), .ZN(n796) );
  NAND2_X1 U891 ( .A1(G104), .A2(n888), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G116), .A2(n883), .ZN(n799) );
  NAND2_X1 U895 ( .A1(G128), .A2(n881), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U897 ( .A(KEYINPUT35), .B(n800), .Z(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U899 ( .A(KEYINPUT36), .B(n803), .ZN(n863) );
  NOR2_X1 U900 ( .A1(n812), .A2(n863), .ZN(n997) );
  NAND2_X1 U901 ( .A1(n997), .A2(n814), .ZN(n809) );
  INV_X1 U902 ( .A(n804), .ZN(n807) );
  XOR2_X1 U903 ( .A(G1986), .B(G290), .Z(n935) );
  NAND2_X1 U904 ( .A1(n1004), .A2(n935), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n805), .A2(n814), .ZN(n806) );
  OR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n816) );
  AND2_X1 U909 ( .A1(n863), .A2(n812), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT104), .ZN(n1015) );
  NAND2_X1 U911 ( .A1(n1015), .A2(n814), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n818) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n817) );
  XNOR2_X1 U914 ( .A(n818), .B(n817), .ZN(G329) );
  XNOR2_X1 U915 ( .A(G2427), .B(G2443), .ZN(n828) );
  XOR2_X1 U916 ( .A(G2430), .B(KEYINPUT107), .Z(n820) );
  XNOR2_X1 U917 ( .A(G2454), .B(G2435), .ZN(n819) );
  XNOR2_X1 U918 ( .A(n820), .B(n819), .ZN(n824) );
  XOR2_X1 U919 ( .A(G2438), .B(KEYINPUT106), .Z(n822) );
  XNOR2_X1 U920 ( .A(G1348), .B(G1341), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U922 ( .A(n824), .B(n823), .Z(n826) );
  XNOR2_X1 U923 ( .A(G2446), .B(G2451), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n829), .A2(G14), .ZN(n905) );
  XOR2_X1 U927 ( .A(KEYINPUT108), .B(n905), .Z(G401) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U930 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n836), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n838) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U943 ( .A(G2678), .B(G2090), .Z(n840) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U945 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U946 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1986), .B(G1971), .Z(n846) );
  XNOR2_X1 U950 ( .A(G1956), .B(G1966), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1976), .Z(n851) );
  XNOR2_X1 U956 ( .A(G1961), .B(G1981), .ZN(n850) );
  XNOR2_X1 U957 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U958 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n881), .ZN(n854) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n854), .Z(n855) );
  XNOR2_X1 U961 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U962 ( .A1(G112), .A2(n883), .ZN(n856) );
  NAND2_X1 U963 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G136), .A2(n516), .ZN(n859) );
  NAND2_X1 U965 ( .A1(G100), .A2(n888), .ZN(n858) );
  NAND2_X1 U966 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U967 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U968 ( .A(n863), .B(n862), .Z(n871) );
  NAND2_X1 U969 ( .A1(G139), .A2(n516), .ZN(n865) );
  NAND2_X1 U970 ( .A1(G103), .A2(n888), .ZN(n864) );
  NAND2_X1 U971 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G115), .A2(n883), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G127), .A2(n881), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n1005) );
  XNOR2_X1 U977 ( .A(n871), .B(n1005), .ZN(n875) );
  XOR2_X1 U978 ( .A(G160), .B(n872), .Z(n873) );
  XNOR2_X1 U979 ( .A(n873), .B(n998), .ZN(n874) );
  XOR2_X1 U980 ( .A(n875), .B(n874), .Z(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n877) );
  XNOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n876) );
  XNOR2_X1 U983 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U984 ( .A(KEYINPUT46), .B(n878), .ZN(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n897) );
  NAND2_X1 U986 ( .A1(n881), .A2(G130), .ZN(n882) );
  XNOR2_X1 U987 ( .A(n882), .B(KEYINPUT110), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n886), .B(KEYINPUT111), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G142), .A2(n516), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n894), .B(G162), .ZN(n895) );
  XOR2_X1 U997 ( .A(G164), .B(n895), .Z(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U999 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(n899), .Z(G395) );
  XNOR2_X1 U1001 ( .A(n949), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(G171), .B(n943), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n903), .B(G286), .ZN(n904) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n904), .ZN(G397) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n905), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1009 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1014 ( .A(G2084), .B(KEYINPUT54), .Z(n911) );
  XNOR2_X1 U1015 ( .A(G34), .B(n911), .ZN(n928) );
  XNOR2_X1 U1016 ( .A(G2090), .B(G35), .ZN(n926) );
  XNOR2_X1 U1017 ( .A(G32), .B(n912), .ZN(n913) );
  NAND2_X1 U1018 ( .A1(n913), .A2(G28), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(G2067), .B(G26), .ZN(n915) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n914) );
  NOR2_X1 U1021 ( .A1(n915), .A2(n914), .ZN(n921) );
  XOR2_X1 U1022 ( .A(n916), .B(G27), .Z(n919) );
  XOR2_X1 U1023 ( .A(n917), .B(G25), .Z(n918) );
  NOR2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n924), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT120), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT55), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(G29), .A2(n931), .ZN(n989) );
  XNOR2_X1 U1033 ( .A(G16), .B(KEYINPUT56), .ZN(n958) );
  XNOR2_X1 U1034 ( .A(n932), .B(G1956), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(n933), .B(KEYINPUT122), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(G166), .B(G1971), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT123), .ZN(n942) );
  XOR2_X1 U1041 ( .A(G171), .B(G1961), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n946) );
  XOR2_X1 U1043 ( .A(G1348), .B(n943), .Z(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(n944), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(n949), .B(G1341), .ZN(n954) );
  XOR2_X1 U1048 ( .A(G168), .B(G1966), .Z(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(KEYINPUT57), .B(n952), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n987) );
  INV_X1 U1054 ( .A(G16), .ZN(n985) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n961) );
  XOR2_X1 U1056 ( .A(G23), .B(KEYINPUT126), .Z(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(G1976), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1059 ( .A(KEYINPUT125), .B(G1971), .Z(n962) );
  XNOR2_X1 U1060 ( .A(G22), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(n965), .Z(n982) );
  XNOR2_X1 U1063 ( .A(G20), .B(n966), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n971) );
  XNOR2_X1 U1069 ( .A(G4), .B(n971), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(KEYINPUT60), .B(n974), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n975), .B(G5), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1076 ( .A(KEYINPUT124), .B(n980), .Z(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n983), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n990), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(KEYINPUT127), .ZN(n1021) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT117), .B(n994), .Z(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT51), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1013) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT116), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G2072), .B(n1005), .Z(n1007) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT118), .B(n1008), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .Z(n1017) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT119), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(G29), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

