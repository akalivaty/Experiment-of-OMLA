//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n209), .A3(new_n206), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT14), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT89), .B(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(G36gat), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n212), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(new_n214), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n211), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n224), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(new_n216), .B2(KEYINPUT15), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n226), .B1(new_n232), .B2(new_n223), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT90), .B1(new_n233), .B2(KEYINPUT17), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT91), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n211), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n211), .A2(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n228), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n233), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n243), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n238), .B(KEYINPUT13), .Z(new_n249));
  AOI22_X1  g048(.A1(new_n244), .A2(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT11), .B(G169gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT12), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n238), .A4(new_n243), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n250), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n250), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n202), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(new_n249), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n257), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n255), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n256), .A3(new_n257), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(KEYINPUT92), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272));
  INV_X1    g071(.A(G211gat), .ZN(new_n273));
  INV_X1    g072(.A(G218gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G211gat), .B(G218gat), .Z(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT72), .ZN(new_n283));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(KEYINPUT24), .A3(new_n287), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n294), .A4(new_n292), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n302), .A2(KEYINPUT28), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n291), .B1(new_n306), .B2(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(KEYINPUT26), .B2(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n283), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n283), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n299), .B2(new_n309), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n281), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n283), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n280), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n318), .A2(new_n319), .A3(new_n314), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n270), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  OR3_X1    g120(.A1(new_n318), .A2(new_n319), .A3(new_n314), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n315), .A3(KEYINPUT74), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(KEYINPUT37), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  NOR2_X1   g126(.A1(new_n316), .A2(new_n320), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n269), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(G141gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n337), .B2(KEYINPUT2), .ZN(new_n338));
  INV_X1    g137(.A(new_n332), .ZN(new_n339));
  INV_X1    g138(.A(G148gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  INV_X1    g141(.A(G141gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(G148gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n333), .B(new_n338), .C1(new_n341), .C2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G141gat), .B(G148gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n334), .B(new_n337), .C1(new_n346), .C2(KEYINPUT2), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(G120gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT1), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n352), .B2(new_n353), .ZN(new_n355));
  OR2_X1    g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356));
  INV_X1    g155(.A(G134gat), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT65), .B(G127gat), .Z(new_n358));
  OAI211_X1 g157(.A(new_n355), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G127gat), .B(G134gat), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT66), .B(G120gat), .Z(new_n361));
  OAI211_X1 g160(.A(new_n354), .B(new_n360), .C1(new_n361), .C2(new_n352), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n363), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n364), .A2(KEYINPUT5), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n345), .A2(new_n350), .A3(new_n369), .A4(new_n349), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n370), .A2(new_n363), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n351), .A2(new_n372), .A3(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n379), .A3(new_n362), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n379), .B1(new_n359), .B2(new_n362), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n347), .B(new_n348), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n333), .A2(new_n338), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n344), .B1(new_n332), .B2(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n345), .A2(new_n350), .A3(KEYINPUT81), .A4(new_n349), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n383), .A2(new_n389), .A3(KEYINPUT4), .A4(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n378), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n365), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n383), .A2(new_n389), .A3(new_n377), .A4(new_n390), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT4), .B1(new_n351), .B2(new_n363), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT5), .B1(new_n396), .B2(new_n375), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n368), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT80), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n351), .A2(new_n372), .A3(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n408), .A2(new_n371), .B1(new_n394), .B2(new_n395), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n392), .B(new_n365), .C1(new_n409), .C2(KEYINPUT5), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n402), .A3(new_n368), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n403), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n269), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n312), .A2(new_n281), .A3(new_n314), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n319), .B1(new_n318), .B2(new_n314), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(KEYINPUT37), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n330), .A2(new_n420), .B1(new_n328), .B2(new_n327), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n415), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n331), .B1(new_n422), .B2(KEYINPUT87), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n402), .B(new_n412), .C1(new_n410), .C2(new_n368), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n414), .B1(new_n398), .B2(new_n403), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n411), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n421), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(G106gat), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n278), .B2(new_n279), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n369), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n278), .C2(new_n279), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n351), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n281), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n370), .A2(new_n311), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n437), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n438), .B(KEYINPUT83), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT3), .B1(new_n280), .B2(new_n311), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n389), .B2(new_n390), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n280), .B1(new_n370), .B2(new_n311), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n442), .B2(new_n447), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n450), .A2(G78gat), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G78gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n442), .A2(new_n447), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G22gat), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n455), .B2(new_n449), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n432), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(G78gat), .B1(new_n450), .B2(new_n451), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n453), .A3(new_n449), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n431), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n396), .A2(new_n375), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n366), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n466), .A2(KEYINPUT85), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(KEYINPUT39), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n402), .B1(new_n465), .B2(KEYINPUT39), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n469), .A3(KEYINPUT40), .ZN(new_n474));
  INV_X1    g273(.A(new_n327), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n321), .A2(new_n475), .A3(new_n323), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n328), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n322), .A2(new_n315), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n475), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n472), .A2(new_n474), .A3(new_n404), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n429), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n381), .B2(new_n382), .ZN(new_n488));
  INV_X1    g287(.A(new_n382), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT68), .A3(new_n380), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n490), .A3(new_n310), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n380), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n492), .A2(new_n487), .A3(new_n299), .A4(new_n309), .ZN(new_n493));
  INV_X1    g292(.A(G227gat), .ZN(new_n494));
  INV_X1    g293(.A(G233gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G15gat), .B(G43gat), .Z(new_n501));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n497), .B(KEYINPUT32), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n493), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT34), .B1(new_n509), .B2(new_n496), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(new_n511), .C1(new_n494), .C2(new_n495), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n504), .A2(new_n510), .A3(new_n512), .A4(new_n506), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n504), .A2(new_n506), .B1(new_n510), .B2(new_n512), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n507), .A2(KEYINPUT69), .A3(new_n513), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n521), .A2(KEYINPUT36), .A3(new_n522), .A4(new_n515), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n524), .A3(new_n517), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n476), .A2(new_n477), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n476), .B2(new_n477), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n481), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n461), .B1(new_n426), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n486), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n534), .A2(new_n457), .A3(new_n460), .ZN(new_n535));
  INV_X1    g334(.A(new_n426), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n515), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n535), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n515), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n461), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n426), .A2(new_n530), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n268), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT94), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n551), .B2(KEYINPUT7), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT95), .A3(G85gat), .A4(G92gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n558), .A3(KEYINPUT7), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n553), .A2(new_n555), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT8), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(G99gat), .B2(G106gat), .ZN(new_n564));
  AND2_X1   g363(.A1(KEYINPUT96), .A2(G92gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(KEYINPUT96), .A2(G92gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n560), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n562), .B1(new_n560), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n228), .B2(new_n229), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n235), .B2(new_n236), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n228), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n453), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n590), .C1(new_n587), .C2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G127gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n246), .B1(new_n598), .B2(new_n597), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT93), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n335), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n605), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n597), .B1(new_n570), .B2(new_n571), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n560), .A2(new_n569), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n561), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n595), .A2(new_n596), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n560), .A2(new_n562), .A3(new_n569), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n622), .A3(KEYINPUT97), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n572), .A2(new_n626), .A3(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n627), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n632), .B2(new_n629), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n634), .B(KEYINPUT10), .C1(new_n623), .C2(new_n627), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n624), .B(KEYINPUT100), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n628), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n643), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n628), .B(new_n645), .C1(new_n637), .C2(new_n625), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n586), .A2(new_n616), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n550), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n426), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n482), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n655), .A2(KEYINPUT101), .B1(KEYINPUT42), .B2(new_n209), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT101), .B2(new_n655), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n658), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n655), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n651), .B2(new_n526), .ZN(new_n665));
  INV_X1    g464(.A(new_n540), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n651), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n462), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND3_X1  g470(.A1(new_n533), .A2(new_n549), .A3(KEYINPUT105), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n484), .B1(new_n423), .B2(new_n428), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n526), .A2(new_n531), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT35), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n545), .B2(new_n546), .ZN(new_n676));
  OAI22_X1  g475(.A1(new_n673), .A2(new_n674), .B1(new_n676), .B2(new_n541), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n586), .A2(KEYINPUT44), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n672), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n586), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n647), .B(KEYINPUT103), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n265), .A2(new_n266), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n615), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT104), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n685), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n215), .B1(new_n694), .B2(new_n536), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n586), .A2(new_n616), .A3(new_n647), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n550), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(new_n536), .A3(new_n215), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(G1328gat));
  INV_X1    g499(.A(new_n482), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n550), .A2(new_n220), .A3(new_n482), .A4(new_n696), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n702), .B(new_n707), .C1(new_n705), .C2(new_n703), .ZN(G1329gat));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n550), .A2(new_n709), .A3(new_n540), .A4(new_n696), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n690), .A2(new_n526), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT47), .B(new_n710), .C1(new_n711), .C2(new_n709), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g514(.A(new_n710), .ZN(new_n716));
  INV_X1    g515(.A(new_n526), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n691), .A2(new_n717), .A3(new_n693), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(G43gat), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n714), .A2(new_n715), .B1(KEYINPUT47), .B2(new_n719), .ZN(G1330gat));
  OAI21_X1  g519(.A(G50gat), .B1(new_n690), .B2(new_n462), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n697), .A2(G50gat), .A3(new_n462), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n691), .A2(new_n461), .A3(new_n693), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n722), .B1(new_n725), .B2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n672), .A2(new_n679), .ZN(new_n728));
  NOR4_X1   g527(.A1(new_n686), .A2(new_n687), .A3(new_n615), .A4(new_n682), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n536), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT109), .B(G57gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n701), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n730), .B2(new_n526), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n540), .A2(new_n589), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g541(.A1(new_n730), .A2(new_n462), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n453), .ZN(G1335gat));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n677), .A2(KEYINPUT110), .A3(new_n682), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n687), .A2(new_n616), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT110), .B1(new_n677), .B2(new_n682), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n683), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n747), .A4(new_n746), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n648), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n568), .A3(new_n426), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n747), .A2(new_n647), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n685), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n536), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(G1336gat));
  NOR2_X1   g559(.A1(new_n701), .A2(G92gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n686), .B(new_n762), .C1(new_n750), .C2(new_n753), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n681), .B2(new_n684), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n567), .B1(new_n764), .B2(new_n482), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(new_n567), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n758), .B2(new_n701), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n769), .B2(KEYINPUT111), .ZN(new_n770));
  INV_X1    g569(.A(new_n686), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n746), .A2(new_n747), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT51), .B1(new_n772), .B2(new_n752), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n748), .A2(new_n745), .A3(new_n749), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n771), .B(new_n761), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n769), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n766), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n770), .B1(new_n766), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n754), .A2(new_n781), .A3(new_n540), .ZN(new_n782));
  OAI21_X1  g581(.A(G99gat), .B1(new_n758), .B2(new_n526), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1338gat));
  NOR2_X1   g583(.A1(new_n462), .A2(G106gat), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n771), .B(new_n785), .C1(new_n773), .C2(new_n774), .ZN(new_n786));
  OAI21_X1  g585(.A(G106gat), .B1(new_n758), .B2(new_n462), .ZN(new_n787));
  NAND2_X1  g586(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n789), .B(new_n790), .Z(G1339gat));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n632), .A2(new_n629), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n634), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n632), .A2(KEYINPUT98), .A3(new_n629), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n625), .B1(new_n796), .B2(new_n631), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n631), .B(new_n638), .C1(new_n633), .C2(new_n635), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT54), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT55), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  INV_X1    g600(.A(new_n638), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n636), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n643), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n646), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n643), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT54), .B(new_n798), .C1(new_n637), .C2(new_n625), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n792), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n797), .A2(new_n799), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n804), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n643), .A4(new_n803), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT114), .A4(new_n646), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n687), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n238), .B1(new_n237), .B2(new_n243), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n248), .A2(new_n249), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n254), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n266), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n648), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n586), .A3(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n809), .A2(new_n814), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n586), .A2(new_n819), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n616), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n649), .A2(new_n687), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n461), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n536), .A2(new_n482), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n666), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n352), .A3(new_n268), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n832), .A2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n545), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n687), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n352), .B2(new_n842), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n361), .A3(new_n647), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n833), .A2(new_n771), .A3(new_n836), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(G120gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(G120gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(G1341gat));
  NAND3_X1  g648(.A1(new_n841), .A2(new_n358), .A3(new_n616), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n837), .A2(new_n615), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n358), .B2(new_n851), .ZN(G1342gat));
  NAND2_X1  g651(.A1(new_n682), .A2(new_n357), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n840), .A2(KEYINPUT56), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n837), .B2(new_n586), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT56), .B1(new_n840), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n717), .A2(new_n462), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n268), .A2(G141gat), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n839), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n717), .A2(new_n835), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n832), .B2(new_n462), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n462), .A2(new_n863), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n268), .A2(new_n805), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n811), .A2(new_n804), .A3(KEYINPUT117), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT117), .B1(new_n811), .B2(new_n804), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n810), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n820), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n829), .B1(new_n870), .B2(new_n682), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n615), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n865), .B1(new_n872), .B2(new_n831), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n862), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n687), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n860), .B1(new_n875), .B2(new_n339), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  INV_X1    g676(.A(new_n268), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n332), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n860), .A2(KEYINPUT58), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n876), .A2(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n648), .A2(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n839), .A2(new_n858), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT118), .Z(new_n884));
  AOI211_X1 g683(.A(KEYINPUT59), .B(new_n340), .C1(new_n874), .C2(new_n647), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n861), .A2(new_n647), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n865), .B1(new_n830), .B2(new_n831), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n878), .A2(new_n649), .A3(KEYINPUT119), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT119), .B1(new_n878), .B2(new_n649), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n828), .A2(new_n646), .A3(new_n813), .A4(new_n812), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n870), .B2(new_n682), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n893), .B2(new_n615), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n863), .B1(new_n894), .B2(new_n462), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n887), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n340), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n886), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n884), .B1(new_n885), .B2(new_n899), .ZN(G1345gat));
  NAND2_X1  g699(.A1(new_n839), .A2(new_n858), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(KEYINPUT121), .A3(new_n615), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(G155gat), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n901), .B2(new_n615), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n615), .A2(new_n335), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n903), .A2(new_n904), .B1(new_n874), .B2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n874), .A2(G162gat), .A3(new_n682), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n336), .B1(new_n901), .B2(new_n586), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NAND3_X1  g708(.A1(new_n540), .A2(new_n536), .A3(new_n482), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n833), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n289), .A3(new_n268), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n830), .A2(new_n831), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n426), .A2(new_n701), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(new_n545), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n687), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n913), .A2(new_n917), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n912), .B2(new_n686), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n290), .A3(new_n647), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1349gat));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n616), .A2(new_n300), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n914), .A2(new_n462), .A3(new_n616), .A4(new_n911), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G183gat), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n923), .B(new_n924), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n922), .A2(new_n926), .A3(new_n928), .A4(KEYINPUT60), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n912), .B2(new_n586), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n301), .A3(new_n682), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n934), .B(new_n935), .C1(new_n938), .C2(new_n939), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n888), .A2(new_n895), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n526), .A2(new_n915), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n268), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n832), .A2(new_n462), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n943), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G197gat), .B1(new_n265), .B2(new_n266), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n948), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  OAI21_X1  g751(.A(G204gat), .B1(new_n944), .B2(new_n686), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n648), .A2(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n946), .A2(new_n943), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT62), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(KEYINPUT62), .ZN(new_n958));
  OAI221_X1 g757(.A(new_n953), .B1(KEYINPUT62), .B2(new_n955), .C1(new_n957), .C2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n948), .A2(new_n273), .A3(new_n616), .ZN(new_n960));
  AOI211_X1 g759(.A(new_n615), .B(new_n942), .C1(new_n888), .C2(new_n895), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n273), .B1(new_n961), .B2(KEYINPUT127), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n942), .B1(new_n888), .B2(new_n895), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT127), .B1(new_n963), .B2(new_n616), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n941), .A2(KEYINPUT127), .A3(new_n616), .A4(new_n943), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G211gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n968), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n960), .B1(new_n966), .B2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n944), .B2(new_n586), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n682), .A2(new_n274), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n947), .B2(new_n973), .ZN(G1355gat));
endmodule


