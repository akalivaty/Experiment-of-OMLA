//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G64gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  OR2_X1    g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT9), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212));
  AOI22_X1  g011(.A1(new_n204), .A2(new_n208), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT21), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n214), .B(new_n215), .Z(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT16), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n222), .A2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  AOI21_X1  g026(.A(G8gat), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(KEYINPUT93), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n213), .A2(KEYINPUT93), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT21), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(G231gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n238), .A2(new_n239), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G155gat), .ZN(new_n243));
  INV_X1    g042(.A(G211gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n238), .A2(new_n239), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n217), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n245), .B1(new_n241), .B2(new_n242), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n248), .A2(new_n240), .A3(new_n247), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n216), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  AND3_X1   g054(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n256));
  XOR2_X1   g055(.A(G43gat), .B(G50gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT14), .Z(new_n261));
  XOR2_X1   g060(.A(KEYINPUT86), .B(G29gat), .Z(new_n262));
  AND3_X1   g061(.A1(new_n262), .A2(KEYINPUT87), .A3(G36gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT87), .B1(new_n262), .B2(G36gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n259), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n257), .A2(new_n258), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  INV_X1    g069(.A(G85gat), .ZN(new_n271));
  INV_X1    g070(.A(G92gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(KEYINPUT8), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT7), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n271), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G99gat), .B(G106gat), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n277), .B(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n256), .B1(new_n269), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n265), .A2(new_n266), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n265), .A2(new_n266), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n267), .A2(KEYINPUT17), .A3(new_n268), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n281), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT94), .ZN(new_n289));
  XOR2_X1   g088(.A(G190gat), .B(G218gat), .Z(new_n290));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n281), .B(new_n291), .C1(new_n287), .C2(new_n280), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n255), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(KEYINPUT95), .A3(new_n293), .ZN(new_n298));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n298), .A3(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n255), .B(new_n301), .C1(new_n294), .C2(new_n295), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n254), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n278), .A2(KEYINPUT96), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n280), .A2(new_n213), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n213), .A2(new_n307), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n277), .B(new_n278), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT10), .B(new_n280), .C1(new_n233), .C2(new_n234), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT10), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n308), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI211_X1 g121(.A(KEYINPUT97), .B(new_n314), .C1(new_n317), .C2(new_n319), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G176gat), .B(G204gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT98), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(G120gat), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(KEYINPUT99), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT99), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n320), .A2(new_n321), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n315), .B1(new_n333), .B2(new_n323), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n320), .B2(new_n316), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n306), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT100), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT100), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n306), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n231), .A2(new_n268), .A3(new_n267), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n269), .A2(new_n229), .A3(new_n230), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G229gat), .A2(G233gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n348), .B(KEYINPUT13), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n285), .A2(new_n231), .A3(new_n286), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT18), .A3(new_n346), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n346), .A3(new_n348), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT18), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT91), .ZN(new_n358));
  XNOR2_X1  g157(.A(G113gat), .B(G141gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G169gat), .B(G197gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n363), .B(KEYINPUT12), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n354), .B(new_n357), .C1(new_n358), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n358), .A3(new_n352), .ZN(new_n367));
  INV_X1    g166(.A(new_n357), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n367), .B(new_n364), .C1(new_n368), .C2(new_n353), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT29), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT24), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n381));
  INV_X1    g180(.A(G190gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n237), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT64), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G169gat), .ZN(new_n387));
  INV_X1    g186(.A(G176gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OR3_X1    g188(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n380), .A2(new_n383), .A3(KEYINPUT64), .A4(new_n381), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n386), .A2(new_n392), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n382), .A2(KEYINPUT66), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G190gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT67), .B1(new_n237), .B2(KEYINPUT27), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT27), .B(G183gat), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(KEYINPUT67), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT28), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n396), .B2(new_n398), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n402), .A2(new_n403), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT26), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(G169gat), .B2(G176gat), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n378), .B(new_n406), .C1(new_n389), .C2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n395), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n399), .A2(new_n237), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n380), .A2(KEYINPUT65), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n380), .A2(new_n381), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(KEYINPUT65), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n393), .B1(new_n414), .B2(new_n392), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n377), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT72), .B(KEYINPUT22), .Z(new_n417));
  NAND2_X1  g216(.A1(G211gat), .A2(G218gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G218gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n244), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n418), .ZN(new_n422));
  XNOR2_X1  g221(.A(G197gat), .B(G204gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n418), .B(new_n421), .C1(new_n425), .C2(new_n417), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n409), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n399), .A2(new_n400), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(G183gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT28), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n404), .A2(new_n401), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT66), .B(G190gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n412), .B1(new_n438), .B2(G183gat), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT65), .B1(new_n380), .B2(new_n381), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n392), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT25), .ZN(new_n442));
  INV_X1    g241(.A(new_n375), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n437), .A2(new_n442), .A3(new_n443), .A4(new_n395), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n416), .A2(new_n427), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n427), .B1(new_n416), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n372), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n416), .A2(new_n444), .ZN(new_n448));
  INV_X1    g247(.A(new_n427), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT73), .ZN(new_n451));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G64gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(new_n272), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n416), .A2(new_n427), .A3(new_n444), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT73), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n446), .A2(new_n372), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT30), .A4(new_n455), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n329), .A2(G141gat), .ZN(new_n465));
  INV_X1    g264(.A(G141gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G148gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT2), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G155gat), .B(G162gat), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G155gat), .ZN(new_n473));
  INV_X1    g272(.A(G162gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n477), .A2(new_n478), .A3(new_n468), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n477), .B2(new_n468), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G127gat), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n482), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G134gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G127gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(G134gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT68), .ZN(new_n488));
  INV_X1    g287(.A(G120gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G113gat), .ZN(new_n490));
  INV_X1    g289(.A(G113gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G120gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT1), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n484), .A2(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n486), .A2(new_n487), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n493), .A2(new_n496), .A3(new_n494), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT4), .B1(new_n481), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n477), .A2(new_n468), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT74), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n477), .A2(new_n478), .A3(new_n468), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT1), .B1(new_n490), .B2(new_n492), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  XNOR2_X1  g305(.A(G127gat), .B(G134gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n483), .B1(new_n507), .B2(KEYINPUT68), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n508), .B2(new_n505), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(new_n504), .A3(new_n509), .A4(new_n472), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(KEYINPUT75), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n481), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n504), .A4(new_n509), .ZN(new_n514));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n481), .A2(KEYINPUT3), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n472), .C1(new_n479), .C2(new_n480), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n498), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n511), .A2(new_n514), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT5), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n481), .B(new_n498), .ZN(new_n522));
  INV_X1    g321(.A(new_n515), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n510), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n526), .A2(new_n519), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G1gat), .B(G29gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G57gat), .B(G85gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT81), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n464), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n519), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n523), .ZN(new_n542));
  AOI211_X1 g341(.A(KEYINPUT82), .B(new_n515), .C1(new_n526), .C2(new_n519), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n522), .A2(new_n523), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(KEYINPUT84), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n546), .A3(KEYINPUT39), .A4(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT39), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n542), .B2(new_n543), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n550), .A2(KEYINPUT83), .A3(new_n536), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT83), .B1(new_n550), .B2(new_n536), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT40), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(KEYINPUT40), .B(new_n548), .C1(new_n551), .C2(new_n552), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT3), .B1(new_n427), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(new_n512), .ZN(new_n560));
  NAND2_X1  g359(.A1(G228gat), .A2(G233gat), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n427), .B1(new_n518), .B2(new_n558), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n424), .A2(KEYINPUT79), .A3(new_n426), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n558), .C1(KEYINPUT79), .C2(new_n424), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n512), .B1(new_n565), .B2(new_n517), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  INV_X1    g366(.A(G22gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G78gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G50gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n563), .A2(new_n567), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G22gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(KEYINPUT80), .A3(new_n569), .A4(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n524), .A2(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n582));
  INV_X1    g381(.A(new_n535), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n535), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n525), .A2(new_n529), .A3(new_n583), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n538), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n585), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n456), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n460), .B2(new_n461), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n447), .A2(new_n451), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n597), .B2(KEYINPUT38), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n455), .A2(KEYINPUT38), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n445), .B2(new_n446), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n596), .A2(new_n600), .A3(new_n454), .A4(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n592), .A2(new_n598), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n557), .A2(new_n581), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n464), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT77), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n606), .A3(new_n589), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n590), .B2(new_n589), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n608), .A2(new_n609), .A3(new_n584), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n585), .A2(new_n588), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n581), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT69), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n498), .B1(new_n410), .B2(new_n415), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n437), .A2(new_n442), .A3(new_n509), .A4(new_n395), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G227gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n374), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  AOI211_X1 g422(.A(KEYINPUT69), .B(new_n623), .C1(new_n617), .C2(new_n618), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT32), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n622), .B2(new_n624), .ZN(new_n627));
  XNOR2_X1  g426(.A(G15gat), .B(G43gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G71gat), .B(G99gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  OAI221_X1 g431(.A(KEYINPUT32), .B1(new_n626), .B2(new_n632), .C1(new_n622), .C2(new_n624), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n623), .A3(new_n618), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  AND3_X1   g435(.A1(new_n631), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n631), .B2(new_n633), .ZN(new_n638));
  OAI211_X1 g437(.A(KEYINPUT71), .B(new_n615), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(new_n633), .ZN(new_n640));
  INV_X1    g439(.A(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n615), .A2(KEYINPUT71), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n615), .A2(KEYINPUT71), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n631), .A2(new_n636), .A3(new_n633), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n604), .A2(new_n614), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n581), .B(new_n605), .C1(new_n637), .C2(new_n638), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n610), .A2(new_n611), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT35), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n642), .A2(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n585), .A2(new_n588), .A3(new_n591), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n605), .A3(new_n581), .A4(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n650), .A2(new_n653), .B1(new_n656), .B2(new_n652), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n371), .B1(new_n648), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n344), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n651), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n464), .ZN(new_n662));
  AND2_X1   g461(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT42), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(G8gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT101), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(G1325gat));
  AOI21_X1  g468(.A(G15gat), .B1(new_n659), .B2(new_n654), .ZN(new_n670));
  INV_X1    g469(.A(new_n647), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n659), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n672), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n659), .A2(new_n613), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  AOI21_X1  g475(.A(new_n305), .B1(new_n648), .B2(new_n657), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n254), .A2(new_n339), .A3(new_n371), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n262), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n651), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n609), .A2(new_n584), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n607), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n585), .A2(new_n588), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n464), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT103), .B1(new_n687), .B2(new_n581), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n612), .A2(new_n689), .A3(new_n613), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n604), .A2(new_n688), .A3(new_n647), .A4(new_n690), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT44), .B(new_n305), .C1(new_n691), .C2(new_n657), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n648), .A2(new_n657), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n303), .A2(new_n304), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n678), .B(KEYINPUT102), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n651), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n683), .B1(new_n701), .B2(new_n681), .ZN(G1328gat));
  OR3_X1    g501(.A1(new_n679), .A2(G36gat), .A3(new_n605), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(KEYINPUT46), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n464), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G36gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(KEYINPUT46), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT104), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(new_n654), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n679), .A2(G43gat), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n699), .A2(new_n671), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n613), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G50gat), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT48), .B1(new_n717), .B2(KEYINPUT106), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n679), .A2(G50gat), .A3(new_n581), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n717), .B(new_n719), .C1(KEYINPUT106), .C2(KEYINPUT48), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1331gat));
  AOI21_X1  g522(.A(new_n370), .B1(new_n691), .B2(new_n657), .ZN(new_n724));
  INV_X1    g523(.A(new_n339), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n306), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n651), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT107), .B(G57gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n727), .A2(new_n605), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  AND2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n732), .B2(new_n733), .ZN(G1333gat));
  NOR3_X1   g535(.A1(new_n727), .A2(G71gat), .A3(new_n711), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n724), .A2(new_n671), .A3(new_n726), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(G71gat), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1334gat));
  NOR2_X1   g540(.A1(new_n727), .A2(new_n581), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT109), .B(G78gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1335gat));
  INV_X1    g543(.A(new_n254), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n691), .A2(new_n657), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n745), .A2(new_n746), .A3(new_n695), .A4(new_n371), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n749), .A2(new_n339), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n651), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n254), .A2(new_n725), .A3(new_n370), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n692), .B2(new_n696), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT110), .B(new_n753), .C1(new_n692), .C2(new_n696), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n728), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n752), .B1(G85gat), .B2(new_n758), .ZN(G1336gat));
  NOR2_X1   g558(.A1(new_n605), .A2(G92gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n749), .A2(new_n339), .A3(new_n750), .A4(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g561(.A(G92gat), .B1(new_n754), .B2(new_n605), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n605), .B1(new_n756), .B2(new_n757), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(new_n272), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n766), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n766), .B2(KEYINPUT52), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(G1337gat));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n770), .A3(new_n654), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n647), .B1(new_n756), .B2(new_n757), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(G1338gat));
  AND2_X1   g572(.A1(new_n756), .A2(new_n757), .ZN(new_n774));
  OAI21_X1  g573(.A(G106gat), .B1(new_n774), .B2(new_n581), .ZN(new_n775));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n776), .A3(new_n613), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  INV_X1    g578(.A(new_n754), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n780), .B2(new_n613), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n779), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n778), .A2(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n354), .A2(new_n365), .A3(new_n357), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n347), .A2(new_n349), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n348), .B1(new_n351), .B2(new_n346), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n363), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n317), .A2(new_n319), .A3(new_n790), .A4(new_n314), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(KEYINPUT54), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n317), .A2(new_n319), .A3(new_n314), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT112), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n794), .C1(new_n333), .C2(new_n323), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n330), .B1(new_n320), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n799), .A2(KEYINPUT55), .B1(new_n331), .B2(new_n336), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n695), .A2(new_n789), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n370), .A3(new_n802), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n339), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n305), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n254), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n306), .A2(new_n339), .A3(new_n370), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n784), .B1(new_n811), .B2(new_n613), .ZN(new_n812));
  INV_X1    g611(.A(new_n810), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n304), .A2(new_n803), .A3(new_n303), .A4(new_n789), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n805), .A2(new_n806), .B1(new_n303), .B2(new_n304), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n745), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .A3(new_n581), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n728), .A2(new_n464), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n812), .A2(new_n818), .A3(new_n654), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n371), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n811), .A2(new_n728), .A3(new_n649), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n491), .A3(new_n370), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n820), .B2(new_n725), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n489), .A3(new_n339), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n822), .B2(new_n254), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n820), .A2(new_n745), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(G127gat), .ZN(G1342gat));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n485), .A3(new_n695), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT56), .Z(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n820), .B2(new_n305), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1343gat));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n671), .B2(new_n581), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n651), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n647), .A2(KEYINPUT118), .A3(new_n613), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n811), .A2(new_n728), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(KEYINPUT119), .A3(new_n839), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n371), .A2(G141gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n605), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n581), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n798), .A2(KEYINPUT114), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n795), .A2(new_n852), .A3(new_n797), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n800), .A2(new_n370), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n806), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(KEYINPUT116), .A3(new_n806), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n305), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n254), .B1(new_n861), .B2(new_n804), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n850), .B1(new_n862), .B2(new_n810), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n817), .A2(new_n613), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n849), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n850), .C1(new_n862), .C2(new_n810), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n819), .A2(new_n647), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n370), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n846), .B2(new_n847), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n838), .A2(G141gat), .A3(new_n371), .A4(new_n840), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n871), .A2(G141gat), .B1(new_n605), .B2(new_n876), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n873), .A2(new_n875), .B1(new_n877), .B2(new_n874), .ZN(G1344gat));
  NAND4_X1  g677(.A1(new_n844), .A2(new_n329), .A3(new_n339), .A4(new_n605), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n341), .A2(new_n343), .A3(new_n370), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n849), .B(new_n613), .C1(new_n881), .C2(new_n862), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n339), .A3(new_n870), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n339), .A3(new_n870), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(new_n880), .A3(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n879), .B1(new_n886), .B2(new_n888), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n869), .A2(new_n254), .A3(new_n870), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G155gat), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n844), .A2(new_n473), .A3(new_n254), .A4(new_n605), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT121), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1346gat));
  AND3_X1   g696(.A1(new_n869), .A2(G162gat), .A3(new_n870), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n844), .A2(new_n695), .A3(new_n605), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n695), .A2(new_n898), .B1(new_n899), .B2(new_n474), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n651), .A2(new_n605), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n581), .A2(new_n817), .A3(new_n654), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n387), .A3(new_n370), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT122), .Z(new_n904));
  NAND4_X1  g703(.A1(new_n812), .A2(new_n818), .A3(new_n654), .A4(new_n901), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n371), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n902), .B2(new_n339), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n905), .A2(new_n725), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n905), .B2(new_n745), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n254), .A3(new_n401), .ZN(new_n912));
  NAND2_X1  g711(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT124), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n914), .B(new_n917), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n695), .A3(new_n399), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n905), .A2(new_n305), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(G190gat), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n920), .B2(G190gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(G1351gat));
  AND2_X1   g724(.A1(new_n647), .A2(new_n901), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n884), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n371), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n817), .A2(new_n613), .A3(new_n926), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT125), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(G197gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n371), .B2(new_n931), .ZN(G1352gat));
  NAND3_X1  g731(.A1(new_n884), .A2(new_n339), .A3(new_n926), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G204gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n929), .A2(G204gat), .A3(new_n725), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT62), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n884), .A2(new_n254), .A3(new_n926), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n254), .A2(new_n244), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n939), .A2(new_n940), .B1(new_n930), .B2(new_n941), .ZN(G1354gat));
  NOR2_X1   g741(.A1(new_n305), .A2(new_n420), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT127), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n420), .B1(new_n930), .B2(new_n305), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(KEYINPUT126), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1355gat));
endmodule


