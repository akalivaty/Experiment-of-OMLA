

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U320 ( .A(n344), .B(n343), .ZN(n345) );
  INV_X1 U321 ( .A(KEYINPUT66), .ZN(n387) );
  XNOR2_X1 U322 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U323 ( .A(n390), .B(n389), .ZN(n392) );
  XNOR2_X1 U324 ( .A(KEYINPUT48), .B(KEYINPUT107), .ZN(n398) );
  XNOR2_X1 U325 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U326 ( .A(KEYINPUT41), .B(n391), .Z(n548) );
  XNOR2_X1 U327 ( .A(KEYINPUT123), .B(n450), .ZN(n581) );
  XOR2_X1 U328 ( .A(n366), .B(n365), .Z(n554) );
  XNOR2_X1 U329 ( .A(n451), .B(G197GAT), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n453), .B(n452), .ZN(G1352GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT23), .B(G204GAT), .Z(n289) );
  XNOR2_X1 U332 ( .A(G22GAT), .B(G218GAT), .ZN(n288) );
  XNOR2_X1 U333 ( .A(n289), .B(n288), .ZN(n304) );
  XOR2_X1 U334 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n291) );
  XNOR2_X1 U335 ( .A(G197GAT), .B(G211GAT), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U337 ( .A(G50GAT), .B(G162GAT), .Z(n364) );
  XOR2_X1 U338 ( .A(n307), .B(n364), .Z(n293) );
  NAND2_X1 U339 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U341 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n295) );
  XNOR2_X1 U342 ( .A(KEYINPUT22), .B(KEYINPUT80), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U344 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U345 ( .A(G155GAT), .B(KEYINPUT2), .Z(n299) );
  XNOR2_X1 U346 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n408) );
  XNOR2_X1 U348 ( .A(G148GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n300), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U350 ( .A(n408), .B(n333), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(n304), .B(n303), .Z(n462) );
  XOR2_X1 U353 ( .A(G169GAT), .B(G8GAT), .Z(n318) );
  XOR2_X1 U354 ( .A(KEYINPUT87), .B(n318), .Z(n306) );
  NAND2_X1 U355 ( .A1(G226GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n313) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n309), .B(G218GAT), .ZN(n352) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G64GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(G176GAT), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n348) );
  XNOR2_X1 U363 ( .A(n352), .B(n348), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U365 ( .A(KEYINPUT78), .B(G183GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT19), .B(n316), .ZN(n440) );
  XOR2_X1 U369 ( .A(n317), .B(n440), .Z(n500) );
  INV_X1 U370 ( .A(n500), .ZN(n515) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n332) );
  XOR2_X1 U373 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n321) );
  XNOR2_X1 U374 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U376 ( .A(G141GAT), .B(G113GAT), .Z(n323) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G50GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U379 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G43GAT), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n353) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(G22GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n328), .B(G15GAT), .ZN(n379) );
  XNOR2_X1 U385 ( .A(n353), .B(n379), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U387 ( .A(n332), .B(n331), .Z(n544) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U389 ( .A(n333), .B(n363), .ZN(n334) );
  AND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n334), .A2(n335), .ZN(n339) );
  INV_X1 U392 ( .A(n334), .ZN(n337) );
  INV_X1 U393 ( .A(n335), .ZN(n336) );
  NAND2_X1 U394 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND2_X1 U395 ( .A1(n339), .A2(n338), .ZN(n340) );
  XOR2_X1 U396 ( .A(n340), .B(KEYINPUT33), .Z(n346) );
  XOR2_X1 U397 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n342) );
  XNOR2_X1 U398 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n341) );
  XOR2_X1 U399 ( .A(n342), .B(n341), .Z(n344) );
  XOR2_X1 U400 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U401 ( .A(n435), .B(KEYINPUT70), .ZN(n343) );
  XNOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n347), .B(KEYINPUT13), .ZN(n371) );
  XNOR2_X1 U404 ( .A(n371), .B(n348), .ZN(n349) );
  XOR2_X1 U405 ( .A(n350), .B(n349), .Z(n391) );
  NAND2_X1 U406 ( .A1(n544), .A2(n548), .ZN(n351) );
  XNOR2_X1 U407 ( .A(KEYINPUT46), .B(n351), .ZN(n385) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n358) );
  XNOR2_X1 U409 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n355) );
  AND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U412 ( .A(n356), .B(KEYINPUT72), .Z(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U414 ( .A(G92GAT), .B(G106GAT), .Z(n360) );
  XNOR2_X1 U415 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n359) );
  XOR2_X1 U416 ( .A(n360), .B(n359), .Z(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  INV_X1 U419 ( .A(n554), .ZN(n569) );
  XOR2_X1 U420 ( .A(G211GAT), .B(KEYINPUT12), .Z(n368) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(G71GAT), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n383) );
  XOR2_X1 U423 ( .A(G78GAT), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U424 ( .A(G127GAT), .B(G155GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U426 ( .A(n371), .B(KEYINPUT73), .Z(n373) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n377) );
  XNOR2_X1 U431 ( .A(G183GAT), .B(KEYINPUT15), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n443) );
  INV_X1 U436 ( .A(n443), .ZN(n577) );
  AND2_X1 U437 ( .A1(n569), .A2(n443), .ZN(n384) );
  AND2_X1 U438 ( .A1(n385), .A2(n384), .ZN(n386) );
  XOR2_X1 U439 ( .A(n386), .B(KEYINPUT47), .Z(n397) );
  XNOR2_X1 U440 ( .A(n554), .B(KEYINPUT36), .ZN(n580) );
  NAND2_X1 U441 ( .A1(n580), .A2(n577), .ZN(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT45), .B(KEYINPUT104), .Z(n388) );
  BUF_X1 U443 ( .A(n391), .Z(n572) );
  NOR2_X1 U444 ( .A1(n392), .A2(n572), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n393), .B(KEYINPUT105), .ZN(n394) );
  NOR2_X1 U446 ( .A1(n544), .A2(n394), .ZN(n395) );
  XNOR2_X1 U447 ( .A(KEYINPUT106), .B(n395), .ZN(n396) );
  NOR2_X1 U448 ( .A1(n397), .A2(n396), .ZN(n399) );
  XNOR2_X1 U449 ( .A(n399), .B(n398), .ZN(n525) );
  NAND2_X1 U450 ( .A1(n515), .A2(n525), .ZN(n401) );
  XOR2_X1 U451 ( .A(KEYINPUT116), .B(KEYINPUT54), .Z(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n423) );
  XOR2_X1 U453 ( .A(KEYINPUT6), .B(KEYINPUT84), .Z(n403) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G120GAT), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U456 ( .A(KEYINPUT83), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U457 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U459 ( .A(n407), .B(n406), .Z(n413) );
  XOR2_X1 U460 ( .A(G162GAT), .B(n408), .Z(n410) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U463 ( .A(G85GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U465 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n415) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U468 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U469 ( .A(KEYINPUT76), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U470 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U472 ( .A(G113GAT), .B(n420), .Z(n439) );
  XNOR2_X1 U473 ( .A(n439), .B(KEYINPUT4), .ZN(n421) );
  XOR2_X1 U474 ( .A(n422), .B(n421), .Z(n513) );
  INV_X1 U475 ( .A(n513), .ZN(n496) );
  NAND2_X1 U476 ( .A1(n423), .A2(n496), .ZN(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT64), .B(n424), .Z(n449) );
  NAND2_X1 U478 ( .A1(n462), .A2(n449), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n425), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U480 ( .A(G176GAT), .B(G99GAT), .Z(n427) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G190GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U483 ( .A(KEYINPUT79), .B(KEYINPUT65), .Z(n429) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(G15GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U486 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT20), .B(KEYINPUT77), .Z(n433) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U493 ( .A(n441), .B(n440), .Z(n526) );
  INV_X1 U494 ( .A(n526), .ZN(n517) );
  NAND2_X1 U495 ( .A1(n442), .A2(n517), .ZN(n568) );
  NOR2_X1 U496 ( .A1(n568), .A2(n443), .ZN(n446) );
  INV_X1 U497 ( .A(G183GAT), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n444), .B(KEYINPUT120), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(G1350GAT) );
  NOR2_X1 U500 ( .A1(n517), .A2(n462), .ZN(n447) );
  XOR2_X1 U501 ( .A(n447), .B(KEYINPUT26), .Z(n541) );
  INV_X1 U502 ( .A(n541), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n449), .A2(n448), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n581), .A2(n544), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n451) );
  INV_X1 U506 ( .A(n544), .ZN(n557) );
  NOR2_X1 U507 ( .A1(n557), .A2(n572), .ZN(n484) );
  XOR2_X1 U508 ( .A(KEYINPUT16), .B(KEYINPUT75), .Z(n455) );
  NAND2_X1 U509 ( .A1(n577), .A2(n569), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n468) );
  NAND2_X1 U511 ( .A1(n515), .A2(n517), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n462), .A2(n456), .ZN(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n500), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U515 ( .A1(n541), .A2(n463), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n460), .A2(n513), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT89), .B(n461), .Z(n467) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT28), .ZN(n504) );
  INV_X1 U520 ( .A(n504), .ZN(n529) );
  NOR2_X1 U521 ( .A1(n463), .A2(n496), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT88), .ZN(n524) );
  NAND2_X1 U523 ( .A1(n526), .A2(n524), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n529), .A2(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n481) );
  NOR2_X1 U526 ( .A1(n468), .A2(n481), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n469), .B(KEYINPUT90), .ZN(n495) );
  NAND2_X1 U528 ( .A1(n484), .A2(n495), .ZN(n478) );
  NOR2_X1 U529 ( .A1(n496), .A2(n478), .ZN(n470) );
  XOR2_X1 U530 ( .A(KEYINPUT34), .B(n470), .Z(n471) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n500), .A2(n478), .ZN(n473) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT91), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(G1325GAT) );
  NOR2_X1 U535 ( .A1(n478), .A2(n526), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT92), .B(KEYINPUT35), .Z(n475) );
  XNOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT93), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n504), .A2(n478), .ZN(n479) );
  XOR2_X1 U541 ( .A(KEYINPUT94), .B(n479), .Z(n480) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n480), .ZN(G1327GAT) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n487) );
  NOR2_X1 U544 ( .A1(n577), .A2(n481), .ZN(n482) );
  NAND2_X1 U545 ( .A1(n580), .A2(n482), .ZN(n483) );
  XNOR2_X1 U546 ( .A(KEYINPUT37), .B(n483), .ZN(n510) );
  NAND2_X1 U547 ( .A1(n484), .A2(n510), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(KEYINPUT38), .ZN(n493) );
  NOR2_X1 U549 ( .A1(n496), .A2(n493), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n493), .A2(n500), .ZN(n489) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(KEYINPUT95), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(G1329GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT96), .ZN(n491) );
  NOR2_X1 U555 ( .A1(n526), .A2(n493), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n492), .Z(G1330GAT) );
  NOR2_X1 U558 ( .A1(n493), .A2(n504), .ZN(n494) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n494), .Z(G1331GAT) );
  INV_X1 U560 ( .A(n548), .ZN(n560) );
  NOR2_X1 U561 ( .A1(n544), .A2(n560), .ZN(n511) );
  NAND2_X1 U562 ( .A1(n511), .A2(n495), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n496), .A2(n505), .ZN(n498) );
  XNOR2_X1 U564 ( .A(KEYINPUT97), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n500), .A2(n505), .ZN(n501) );
  XOR2_X1 U568 ( .A(KEYINPUT98), .B(n501), .Z(n502) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n526), .A2(n505), .ZN(n503) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n509) );
  XOR2_X1 U573 ( .A(KEYINPUT99), .B(KEYINPUT43), .Z(n507) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT100), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT101), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n520), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n520), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT102), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT103), .B(KEYINPUT44), .Z(n522) );
  NAND2_X1 U587 ( .A1(n520), .A2(n529), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n531) );
  NAND2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n542) );
  NOR2_X1 U592 ( .A1(n526), .A2(n542), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(n527), .Z(n528) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n538), .A2(n544), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n534) );
  NAND2_X1 U599 ( .A1(n538), .A2(n548), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NAND2_X1 U602 ( .A1(n538), .A2(n577), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n554), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n546) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(KEYINPUT112), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n544), .A2(n555), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U615 ( .A1(n555), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(G155GAT), .B(KEYINPUT115), .Z(n553) );
  NAND2_X1 U619 ( .A1(n577), .A2(n555), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n568), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n568), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT118), .B(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1351GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT124), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

