//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n204), .B(new_n205), .C1(G183gat), .C2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n210), .A2(KEYINPUT23), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G190gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n202), .A2(KEYINPUT66), .A3(new_n203), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n217), .B(new_n220), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT25), .B1(new_n225), .B2(G169gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(KEYINPUT23), .B2(new_n207), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n217), .B1(new_n234), .B2(new_n220), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n216), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT27), .B1(new_n237), .B2(KEYINPUT68), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(G183gat), .ZN(new_n241));
  INV_X1    g040(.A(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT27), .B(G183gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(G190gat), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n243), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NOR3_X1   g046(.A1(KEYINPUT69), .A2(G169gat), .A3(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n207), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR4_X1   g049(.A1(KEYINPUT69), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n202), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(G113gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n262), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n224), .A3(new_n229), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n253), .B1(new_n276), .B2(new_n216), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n264), .A2(new_n271), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n281), .B(KEYINPUT64), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G15gat), .B(G43gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n282), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n273), .B2(new_n279), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n292), .B2(KEYINPUT33), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n279), .A3(new_n281), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT34), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n282), .A2(KEYINPUT34), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n273), .A2(new_n279), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n290), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(G22gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G228gat), .ZN(new_n307));
  INV_X1    g106(.A(G233gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G197gat), .ZN(new_n311));
  INV_X1    g110(.A(G204gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G211gat), .A2(G218gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n320), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n313), .A2(new_n314), .B1(new_n317), .B2(new_n316), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(G148gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n331), .B2(G141gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n333), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n331), .A2(G141gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n321), .A2(new_n325), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n335), .A2(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n328), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n326), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n348), .A2(KEYINPUT86), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n327), .B2(new_n328), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT86), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n310), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n319), .B2(new_n320), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n322), .A2(new_n323), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n328), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n309), .B1(new_n361), .B2(new_n347), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(new_n349), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT31), .B(G50gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n357), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n363), .B1(new_n355), .B2(new_n354), .ZN(new_n369));
  INV_X1    g168(.A(new_n356), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n309), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n306), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n366), .B1(new_n357), .B2(new_n365), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n364), .A3(new_n368), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n305), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n302), .B1(new_n290), .B2(new_n296), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n303), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n347), .B2(new_n272), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n278), .A2(new_n381), .A3(new_n350), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n264), .A2(new_n271), .A3(KEYINPUT79), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT79), .B1(new_n264), .B2(new_n271), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n351), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n278), .A2(new_n350), .A3(new_n388), .A4(new_n381), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OR3_X1    g191(.A1(new_n390), .A2(KEYINPUT5), .A3(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT82), .ZN(new_n395));
  XOR2_X1   g194(.A(G57gat), .B(G85gat), .Z(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT5), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n347), .B1(new_n385), .B2(new_n386), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n278), .A2(new_n350), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(new_n392), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n382), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n405), .A3(new_n391), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT80), .B1(new_n404), .B2(new_n406), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n393), .B(new_n399), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n403), .A2(new_n392), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n412), .A3(KEYINPUT5), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n404), .A2(KEYINPUT80), .A3(new_n406), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n399), .B1(new_n417), .B2(new_n393), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT85), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n393), .B1(new_n407), .B2(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(new_n399), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(new_n423), .A3(new_n410), .A4(new_n409), .ZN(new_n424));
  INV_X1    g223(.A(new_n410), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n419), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT77), .ZN(new_n428));
  XOR2_X1   g227(.A(G8gat), .B(G36gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT76), .ZN(new_n430));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT74), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n236), .A2(new_n254), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT29), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n236), .B2(new_n254), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n349), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n236), .A2(new_n254), .A3(new_n434), .ZN(new_n441));
  INV_X1    g240(.A(new_n349), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n277), .C2(new_n437), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT75), .B(new_n349), .C1(new_n435), .C2(new_n438), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n432), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n428), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n445), .ZN(new_n450));
  INV_X1    g249(.A(new_n432), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n445), .A3(new_n432), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n446), .A2(KEYINPUT77), .A3(KEYINPUT30), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n449), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n379), .A2(new_n427), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n293), .A2(new_n295), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n293), .A2(new_n295), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n301), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n290), .A2(new_n296), .A3(new_n302), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(KEYINPUT72), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n378), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n390), .A2(KEYINPUT5), .A3(new_n392), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n415), .B2(new_n416), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT89), .B1(new_n468), .B2(new_n399), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n420), .A2(new_n470), .A3(new_n421), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n410), .A3(new_n471), .A4(new_n409), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n426), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n377), .A2(KEYINPUT35), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n466), .A2(new_n473), .A3(new_n456), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n427), .A2(new_n456), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n377), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n390), .A2(new_n392), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT39), .B1(new_n403), .B2(new_n392), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n390), .A2(new_n484), .A3(new_n392), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n399), .ZN(new_n486));
  NOR2_X1   g285(.A1(KEYINPUT88), .A2(KEYINPUT40), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n483), .B2(new_n486), .ZN(new_n489));
  AND4_X1   g288(.A1(new_n469), .A2(new_n488), .A3(new_n471), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n447), .A2(new_n428), .A3(new_n448), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT77), .B1(new_n446), .B2(KEYINPUT30), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n452), .A4(new_n453), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n450), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n432), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n451), .B1(new_n450), .B2(new_n495), .ZN(new_n500));
  INV_X1    g299(.A(new_n439), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n501), .B2(KEYINPUT90), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n439), .A2(new_n503), .A3(new_n443), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT38), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n446), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n472), .A2(new_n499), .A3(new_n506), .A4(new_n426), .ZN(new_n507));
  INV_X1    g306(.A(new_n377), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n494), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n463), .A2(new_n465), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n461), .A2(KEYINPUT36), .A3(new_n462), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n480), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n476), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT101), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n516), .B2(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT101), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G57gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT99), .B1(new_n525), .B2(G64gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT99), .ZN(new_n527));
  INV_X1    g326(.A(G64gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(G57gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(G64gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT100), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT100), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n526), .A2(new_n529), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n524), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n518), .B1(new_n536), .B2(new_n522), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G127gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G183gat), .B(G211gat), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(G1gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  AOI21_X1  g349(.A(G8gat), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n551), .B(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n539), .B2(new_n538), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  INV_X1    g358(.A(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n558), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n545), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n558), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n563), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n546), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(G43gat), .A2(G50gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(G43gat), .A2(G50gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(KEYINPUT92), .A3(new_n571), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(KEYINPUT15), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G29gat), .A2(G36gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n580));
  INV_X1    g379(.A(G29gat), .ZN(new_n581));
  INV_X1    g380(.A(G36gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n578), .A2(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT94), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n584), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT15), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n572), .B2(new_n573), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n589), .A2(new_n590), .A3(new_n575), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n576), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n586), .A2(new_n593), .B1(new_n576), .B2(new_n596), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT17), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(KEYINPUT8), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n603), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n612), .A3(new_n603), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n602), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n608), .A2(new_n603), .A3(new_n612), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n613), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n598), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n623), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n617), .A2(new_n628), .A3(new_n621), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n627), .B1(new_n624), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n538), .A2(new_n616), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n535), .A3(new_n537), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n619), .A2(new_n537), .A3(new_n535), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT10), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n635), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n643), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n639), .A2(new_n641), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT104), .B1(new_n650), .B2(new_n634), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n652), .B(new_n635), .C1(new_n639), .C2(new_n641), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n648), .B1(new_n654), .B2(new_n647), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n569), .A2(new_n633), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n554), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n551), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n598), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n555), .B1(new_n601), .B2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n598), .A2(new_n599), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n657), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT18), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT96), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(KEYINPUT98), .B1(new_n659), .B2(new_n598), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n659), .B2(new_n598), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n555), .A2(KEYINPUT98), .A3(new_n601), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT97), .B(KEYINPUT13), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n657), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n600), .A2(new_n555), .A3(new_n602), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(new_n657), .A3(new_n660), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G197gat), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT11), .B(G169gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n671), .A3(new_n681), .A4(new_n674), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n656), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n515), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n427), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n493), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G8gat), .B1(new_n688), .B2(new_n456), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n693), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n700), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT105), .B1(new_n702), .B2(new_n697), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1325gat));
  AND2_X1   g503(.A1(new_n463), .A2(new_n465), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n688), .A2(G15gat), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n513), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(G15gat), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT106), .Z(G1326gat));
  INV_X1    g509(.A(new_n479), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n688), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n655), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n569), .A2(new_n686), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n515), .A2(new_n632), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n581), .A3(new_n690), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n480), .A2(new_n509), .A3(new_n513), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n473), .A2(new_n456), .A3(new_n474), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n466), .B1(new_n457), .B2(KEYINPUT35), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT107), .B(new_n632), .C1(new_n720), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n515), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n632), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n726), .A3(new_n716), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n427), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n719), .A2(new_n728), .ZN(G1328gat));
  NAND4_X1  g528(.A1(new_n725), .A2(new_n493), .A3(new_n726), .A4(new_n716), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G36gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n456), .A2(G36gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n515), .A2(new_n632), .A3(new_n716), .A4(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n707), .A3(new_n726), .A4(new_n716), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n743), .A3(new_n466), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT47), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n742), .B(new_n744), .C1(new_n746), .C2(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1330gat));
  OAI21_X1  g549(.A(G50gat), .B1(new_n727), .B2(new_n508), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n711), .A2(G50gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n717), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(KEYINPUT48), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n479), .A3(new_n726), .A4(new_n716), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n755), .A2(G50gat), .B1(new_n717), .B2(new_n752), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g556(.A(new_n569), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n758), .A2(new_n685), .A3(new_n632), .A4(new_n655), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n515), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n427), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n525), .ZN(G1332gat));
  OR2_X1    g561(.A1(new_n493), .A2(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n493), .A2(KEYINPUT110), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  NOR3_X1   g569(.A1(new_n760), .A2(G71gat), .A3(new_n705), .ZN(new_n771));
  INV_X1    g570(.A(new_n760), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n707), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(G71gat), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n479), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g576(.A1(new_n427), .A2(G85gat), .A3(new_n655), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n569), .A2(new_n685), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n515), .A2(new_n632), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n515), .A2(KEYINPUT51), .A3(new_n632), .A4(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n569), .A2(new_n685), .A3(new_n655), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n725), .A2(new_n726), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n427), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1336gat));
  OAI21_X1  g590(.A(G92gat), .B1(new_n789), .B2(new_n765), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n765), .A2(G92gat), .A3(new_n655), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n784), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n780), .A2(new_n796), .A3(KEYINPUT51), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT51), .B1(new_n780), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n725), .A2(new_n493), .A3(new_n726), .A4(new_n788), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n799), .A2(new_n793), .B1(G92gat), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n795), .B1(new_n801), .B2(new_n802), .ZN(G1337gat));
  NOR3_X1   g602(.A1(new_n705), .A2(G99gat), .A3(new_n655), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT113), .Z(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n785), .B2(new_n786), .ZN(new_n806));
  OAI21_X1  g605(.A(G99gat), .B1(new_n789), .B2(new_n513), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1338gat));
  OAI21_X1  g607(.A(G106gat), .B1(new_n789), .B2(new_n508), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n508), .A2(G106gat), .A3(new_n655), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT53), .B1(new_n784), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n725), .A2(new_n479), .A3(new_n726), .A4(new_n788), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n799), .A2(new_n810), .B1(G106gat), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(new_n765), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n427), .A3(new_n705), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n651), .A2(new_n653), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n646), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n650), .B2(new_n634), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n639), .A2(new_n635), .A3(new_n641), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n535), .A2(new_n537), .B1(new_n615), .B2(new_n614), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n640), .A2(new_n828), .A3(KEYINPUT10), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n638), .A2(new_n637), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n634), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n652), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n820), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n826), .B1(new_n822), .B2(new_n823), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n647), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(new_n648), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n685), .B(new_n827), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n670), .B1(new_n667), .B2(new_n668), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n657), .B1(new_n672), .B2(new_n660), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n679), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n684), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n655), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n632), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n632), .B(new_n827), .C1(new_n839), .C2(new_n840), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n845), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n758), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n656), .A2(new_n685), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n479), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n818), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n855), .A2(new_n267), .A3(new_n686), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n690), .ZN(new_n858));
  INV_X1    g657(.A(new_n379), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(new_n817), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n685), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(new_n267), .ZN(G1340gat));
  NOR2_X1   g661(.A1(new_n655), .A2(G120gat), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n855), .B2(new_n655), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n258), .A3(new_n569), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n855), .B2(new_n758), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  NAND2_X1  g669(.A1(new_n456), .A2(new_n632), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n858), .A2(G134gat), .A3(new_n859), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n855), .B2(new_n633), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(G1343gat));
  AOI21_X1  g676(.A(new_n508), .B1(new_n851), .B2(new_n853), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n825), .A2(new_n826), .B1(new_n683), .B2(new_n684), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n836), .A2(new_n838), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n846), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n884), .A2(new_n632), .B1(new_n849), .B2(new_n845), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n852), .B1(new_n885), .B2(new_n758), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n711), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n817), .A2(new_n427), .A3(new_n707), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n880), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(G141gat), .B1(new_n889), .B2(new_n686), .ZN(new_n890));
  INV_X1    g689(.A(new_n858), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n707), .A2(new_n508), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT117), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n686), .A2(G141gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n891), .A2(new_n893), .A3(new_n765), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1344gat));
  AOI21_X1  g699(.A(KEYINPUT55), .B1(new_n821), .B2(new_n824), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n632), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n849), .A2(KEYINPUT119), .ZN(new_n907));
  INV_X1    g706(.A(new_n845), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n686), .A2(new_n901), .A3(new_n882), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n633), .B1(new_n910), .B2(new_n846), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n852), .B1(new_n912), .B2(new_n758), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n711), .A2(KEYINPUT57), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n913), .A2(new_n915), .B1(new_n878), .B2(new_n879), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n715), .ZN(new_n917));
  OAI21_X1  g716(.A(G148gat), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT59), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n880), .A2(new_n887), .A3(new_n715), .A4(new_n888), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n331), .A2(KEYINPUT59), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n920), .A2(KEYINPUT118), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT118), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n891), .A2(new_n893), .A3(new_n765), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n925), .A2(G148gat), .A3(new_n655), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n889), .B2(new_n758), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n569), .A2(new_n560), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n925), .B2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n889), .B2(new_n633), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n871), .A2(G162gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n891), .A2(new_n893), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1347gat));
  NAND2_X1  g733(.A1(new_n427), .A2(new_n493), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n705), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT120), .Z(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n854), .ZN(new_n938));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n686), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n765), .A2(new_n690), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n857), .A2(new_n379), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n941), .A2(new_n210), .A3(new_n212), .A4(new_n685), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n938), .B2(new_n655), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n211), .A3(new_n715), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n938), .B2(new_n758), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT122), .B1(new_n948), .B2(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n245), .A3(new_n569), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n947), .B2(new_n950), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n954), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n242), .A3(new_n632), .ZN(new_n956));
  OAI21_X1  g755(.A(G190gat), .B1(new_n938), .B2(new_n633), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NAND3_X1  g759(.A1(new_n904), .A2(new_n632), .A3(new_n908), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n846), .B1(new_n904), .B2(new_n685), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n632), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n852), .B1(new_n963), .B2(new_n758), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT57), .B1(new_n964), .B2(new_n508), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n569), .B1(new_n909), .B2(new_n911), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n914), .B1(new_n966), .B2(new_n852), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n707), .A2(new_n935), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n965), .A2(new_n685), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G197gat), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n857), .A2(new_n940), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n971), .A2(new_n311), .A3(new_n685), .A4(new_n892), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n975), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1352gat));
  NAND4_X1  g776(.A1(new_n965), .A2(new_n715), .A3(new_n967), .A4(new_n968), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n312), .B1(new_n978), .B2(KEYINPUT124), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(KEYINPUT124), .B2(new_n978), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n971), .A2(new_n312), .A3(new_n715), .A4(new_n892), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT62), .Z(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1353gat));
  NOR2_X1   g782(.A1(new_n758), .A2(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n971), .A2(new_n892), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n965), .A2(new_n569), .A3(new_n967), .A4(new_n968), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G211gat), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT63), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT63), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n990), .A3(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n986), .A2(new_n989), .A3(new_n991), .ZN(G1354gat));
  NOR3_X1   g791(.A1(new_n916), .A2(new_n707), .A3(new_n935), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n632), .A2(G218gat), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n971), .A2(new_n632), .A3(new_n892), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n993), .A2(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G1355gat));
endmodule


