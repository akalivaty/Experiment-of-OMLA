//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AND2_X1   g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G20), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n210), .B1(new_n213), .B2(new_n214), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G1), .A3(G13), .ZN(new_n244));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n246));
  AND2_X1   g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G226), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT69), .A2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT69), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n253), .B1(new_n211), .B2(new_n243), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n254), .A3(new_n245), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n244), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(G190), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G58), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT8), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n202), .ZN(new_n286));
  INV_X1    g0086(.A(new_n282), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G1), .B2(new_n277), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n288), .B2(new_n202), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(KEYINPUT9), .B1(new_n291), .B2(KEYINPUT10), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n283), .A2(new_n289), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n268), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n268), .A2(new_n292), .A3(new_n295), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n265), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n293), .B(new_n302), .C1(G169), .C2(new_n265), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  INV_X1    g0106(.A(G238), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n305), .B1(new_n306), .B2(new_n257), .C1(new_n261), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n264), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n247), .A2(G244), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n255), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G20), .A2(G77), .ZN(new_n314));
  INV_X1    g0114(.A(new_n269), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n271), .B2(new_n315), .C1(new_n278), .C2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n282), .B1(new_n260), .B2(new_n285), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT71), .B1(new_n288), .B2(new_n260), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n282), .B1(new_n245), .B2(G20), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT71), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n311), .B1(new_n308), .B2(new_n264), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n313), .B(new_n324), .C1(G169), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n318), .A2(new_n323), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(G190), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(new_n266), .C2(new_n325), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n260), .B2(new_n278), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n332), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT12), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n285), .B2(new_n330), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n284), .A2(KEYINPUT12), .A3(G68), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n288), .A2(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT11), .B1(new_n332), .B2(new_n282), .ZN(new_n338));
  OR3_X1    g0138(.A1(new_n333), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(KEYINPUT69), .A2(G41), .ZN(new_n340));
  NOR2_X1   g0140(.A1(KEYINPUT69), .A2(G41), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(G1), .B1(new_n342), .B2(new_n250), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n254), .B1(new_n247), .B2(G238), .ZN(new_n344));
  INV_X1    g0144(.A(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(G232), .A4(G1698), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(G226), .A4(new_n258), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n264), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n344), .B2(new_n353), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n339), .B1(new_n357), .B2(G190), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT73), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n344), .A2(new_n353), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G190), .A3(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n333), .A2(new_n337), .A3(new_n338), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT73), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n326), .B(new_n329), .C1(new_n360), .C2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G169), .B1(new_n355), .B2(new_n356), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(G169), .C1(new_n355), .C2(new_n356), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(G179), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n365), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n304), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n346), .A2(new_n348), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT7), .A4(new_n277), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n257), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(G20), .B1(new_n346), .B2(new_n348), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n379), .B1(new_n384), .B2(KEYINPUT7), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n274), .A2(new_n330), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n387), .B2(new_n201), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n269), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n378), .A2(KEYINPUT7), .A3(new_n277), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n330), .B1(new_n382), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n395), .B2(new_n390), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n282), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n276), .A2(new_n320), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n284), .B2(new_n276), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n244), .A2(G232), .A3(new_n246), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n255), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n346), .A2(new_n348), .A3(G226), .A4(G1698), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n346), .A2(new_n348), .A3(G223), .A4(new_n258), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n264), .ZN(new_n408));
  INV_X1    g0208(.A(G190), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n255), .A2(new_n402), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n264), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(G200), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n397), .A2(new_n398), .A3(new_n401), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n257), .A2(new_n381), .A3(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT7), .B1(new_n378), .B2(new_n277), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n391), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n287), .B1(new_n420), .B2(new_n393), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n400), .B1(new_n421), .B2(new_n392), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT76), .A3(new_n398), .A4(new_n413), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n396), .A2(new_n282), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n413), .B(new_n401), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n422), .A2(KEYINPUT75), .A3(new_n413), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n412), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n403), .A2(G179), .A3(new_n408), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n397), .A2(new_n401), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n422), .A2(new_n437), .A3(KEYINPUT18), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n377), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n245), .A2(G33), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n287), .A2(new_n284), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G116), .ZN(new_n447));
  INV_X1    g0247(.A(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n285), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(new_n345), .B2(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT78), .B1(G33), .B2(G283), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n280), .A2(new_n281), .B1(G20), .B2(new_n448), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT20), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n456), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n447), .B(new_n449), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n346), .A2(new_n348), .A3(G264), .A4(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n346), .A2(new_n348), .A3(G257), .A4(new_n258), .ZN(new_n461));
  INV_X1    g0261(.A(G303), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n460), .B(new_n461), .C1(new_n462), .C2(new_n257), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n264), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n245), .B(G45), .C1(new_n465), .C2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n340), .B2(new_n341), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n264), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G270), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n249), .A2(new_n251), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n471), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n254), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n464), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n459), .A2(new_n474), .A3(KEYINPUT21), .A4(G169), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n459), .A2(new_n474), .A3(G169), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n459), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(G200), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n469), .A2(G270), .B1(new_n472), .B2(new_n254), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(G190), .A3(new_n464), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n474), .A2(new_n301), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n459), .ZN(new_n485));
  AND4_X1   g0285(.A1(new_n475), .A2(new_n478), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G97), .A2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(G87), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(new_n351), .B2(new_n277), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G97), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n489), .A2(new_n490), .B1(new_n278), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n257), .A2(KEYINPUT79), .A3(new_n277), .A4(G68), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n346), .A2(new_n348), .A3(new_n277), .A4(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT79), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n282), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n316), .A2(new_n285), .ZN(new_n499));
  INV_X1    g0299(.A(new_n316), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n446), .A2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G250), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n250), .B2(G1), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n245), .A2(new_n253), .A3(G45), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n244), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n346), .A2(new_n348), .A3(G238), .A4(new_n258), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n346), .A2(new_n348), .A3(G244), .A4(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(new_n264), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n301), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G169), .B2(new_n512), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(G190), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n266), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n446), .A2(G87), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n498), .A2(new_n499), .A3(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n502), .A2(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n346), .A2(new_n348), .A3(G250), .A4(new_n258), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n257), .A2(KEYINPUT80), .A3(G250), .A4(new_n258), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n346), .A2(new_n348), .A3(G257), .A4(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n264), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n469), .A2(G264), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n301), .A3(new_n473), .A4(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n346), .A2(new_n348), .A3(new_n277), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n257), .A2(new_n535), .A3(new_n277), .A4(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n510), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n277), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n306), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n538), .B1(new_n537), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n282), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT25), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n284), .B2(G107), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n284), .A2(new_n548), .A3(G107), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n446), .A2(G107), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n527), .B1(new_n522), .B2(new_n523), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n473), .B(new_n531), .C1(new_n553), .C2(new_n244), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n547), .A2(new_n552), .B1(new_n434), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n519), .B1(new_n532), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(G200), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n530), .A2(G190), .A3(new_n473), .A4(new_n531), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n547), .A2(new_n557), .A3(new_n558), .A4(new_n552), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n284), .A2(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n446), .B2(G97), .ZN(new_n561));
  OAI21_X1  g0361(.A(G107), .B1(new_n417), .B2(new_n418), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT6), .ZN(new_n563));
  AND2_X1   g0363(.A1(G97), .A2(G107), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n487), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT6), .A2(G97), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT77), .B1(new_n566), .B2(G107), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT77), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(new_n306), .A3(KEYINPUT6), .A4(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n561), .B1(new_n572), .B2(new_n287), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT5), .B1(new_n249), .B2(new_n251), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n244), .C1(new_n574), .C2(new_n466), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n473), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n346), .A2(new_n348), .A3(G244), .A4(new_n258), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n453), .A2(new_n454), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n576), .B1(new_n264), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n301), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n473), .A2(new_n575), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n264), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n434), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n573), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(G190), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(G200), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n287), .B1(new_n562), .B2(new_n571), .ZN(new_n593));
  INV_X1    g0393(.A(new_n561), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n559), .A2(new_n590), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n444), .A2(new_n486), .A3(new_n556), .A4(new_n597), .ZN(G372));
  OAI22_X1  g0398(.A1(new_n584), .A2(G169), .B1(new_n593), .B2(new_n594), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n588), .A2(G179), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT82), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT82), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n573), .A2(new_n585), .A3(new_n589), .A4(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT26), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n502), .A2(new_n514), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT81), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n518), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n498), .A2(KEYINPUT81), .A3(new_n499), .A4(new_n517), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n516), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n604), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n519), .A2(new_n590), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n606), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n590), .A2(new_n596), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n554), .A2(new_n434), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n537), .A2(new_n543), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT24), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n287), .B1(new_n620), .B2(new_n544), .ZN(new_n621));
  INV_X1    g0421(.A(new_n552), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n532), .B(new_n618), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n476), .A2(new_n477), .B1(new_n484), .B2(new_n459), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n475), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n617), .A2(new_n625), .A3(new_n559), .A4(new_n612), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n613), .A2(new_n615), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n444), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n628), .B(KEYINPUT83), .Z(new_n629));
  INV_X1    g0429(.A(new_n303), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n326), .A2(KEYINPUT84), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n325), .A2(G169), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT84), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n313), .A4(new_n324), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n366), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n432), .B1(new_n376), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n442), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n298), .A2(new_n300), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n629), .A2(new_n641), .ZN(G369));
  NAND3_X1  g0442(.A1(new_n245), .A2(new_n277), .A3(G13), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n459), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n486), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n624), .A2(new_n475), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n623), .A2(new_n648), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n648), .B1(new_n621), .B2(new_n622), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n559), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n623), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n652), .A2(new_n648), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n655), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n612), .A2(KEYINPUT26), .A3(new_n601), .A4(new_n603), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n605), .B1(new_n519), .B2(new_n590), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT87), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n604), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n612), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n652), .A2(new_n671), .A3(new_n623), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n590), .A2(new_n596), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n590), .B2(new_n596), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n612), .A2(new_n559), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n625), .A2(KEYINPUT88), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n672), .A2(new_n676), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n606), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n670), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n648), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n664), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n627), .A2(new_n682), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n530), .A2(new_n531), .A3(new_n587), .A4(new_n586), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n481), .A2(new_n512), .A3(G179), .A4(new_n464), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n690), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n529), .A2(new_n264), .B1(G264), .B2(new_n469), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(KEYINPUT30), .A3(new_n693), .A4(new_n584), .ZN(new_n694));
  AOI21_X1  g0494(.A(G179), .B1(new_n481), .B2(new_n464), .ZN(new_n695));
  INV_X1    g0495(.A(new_n512), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n588), .A2(new_n695), .A3(new_n554), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT31), .B1(new_n698), .B2(new_n648), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n687), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n648), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(KEYINPUT86), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n597), .A2(new_n556), .A3(new_n486), .A4(new_n682), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n701), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n686), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n245), .ZN(new_n711));
  INV_X1    g0511(.A(new_n208), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n471), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G1), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n487), .A2(new_n488), .A3(new_n448), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT85), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n715), .A2(new_n717), .B1(new_n214), .B2(new_n714), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(G364));
  AND2_X1   g0520(.A1(new_n277), .A2(G13), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n245), .B1(new_n721), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OR3_X1    g0523(.A1(new_n723), .A2(new_n713), .A3(KEYINPUT90), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT90), .B1(new_n723), .B2(new_n713), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n654), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n653), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n257), .A2(G355), .A3(new_n208), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G116), .B2(new_n208), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n378), .A2(new_n208), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n214), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(new_n250), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n241), .A2(new_n250), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n281), .B1(G20), .B2(new_n434), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n727), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n277), .A2(G190), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT92), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT92), .ZN(new_n748));
  AND4_X1   g0548(.A1(new_n301), .A2(new_n747), .A3(G200), .A4(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G283), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n747), .A2(new_n748), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT94), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT94), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G329), .ZN(new_n760));
  INV_X1    g0560(.A(new_n746), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n301), .A3(new_n266), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n277), .A2(new_n409), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n301), .A3(G200), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n764), .B1(new_n766), .B2(new_n462), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n761), .A2(new_n301), .A3(G200), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n257), .B(new_n767), .C1(G311), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n765), .A2(G179), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G326), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n765), .A2(G179), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n277), .B1(new_n754), .B2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(G294), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n753), .A2(new_n760), .A3(new_n769), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n752), .A2(G107), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n771), .A2(G50), .B1(new_n779), .B2(G97), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n274), .B2(new_n775), .ZN(new_n784));
  INV_X1    g0584(.A(new_n768), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n257), .B1(new_n785), .B2(new_n260), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n763), .A2(new_n330), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n766), .A2(new_n488), .ZN(new_n788));
  NOR4_X1   g0588(.A1(new_n784), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n755), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n782), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n745), .B1(new_n794), .B2(new_n742), .ZN(new_n795));
  INV_X1    g0595(.A(new_n741), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n653), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n729), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NOR2_X1   g0599(.A1(new_n742), .A2(new_n739), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n727), .B1(G77), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT34), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G150), .A2(new_n762), .B1(new_n768), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT96), .B(G143), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n770), .C1(new_n775), .C2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n803), .A2(new_n807), .B1(new_n759), .B2(G132), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n378), .B1(new_n779), .B2(G58), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(new_n803), .C2(new_n807), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n752), .A2(G68), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n202), .B2(new_n766), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n812), .B2(KEYINPUT97), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(KEYINPUT97), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n758), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n752), .A2(G87), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n378), .B1(new_n766), .B2(new_n306), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT95), .Z(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n775), .A2(new_n820), .B1(new_n770), .B2(new_n462), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n785), .A2(new_n448), .B1(new_n763), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(G97), .C2(new_n779), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n817), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n814), .B1(new_n816), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n802), .B1(new_n826), .B2(new_n742), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT98), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n324), .A2(new_n648), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n329), .A2(new_n326), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT99), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n329), .A2(KEYINPUT99), .A3(new_n326), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  INV_X1    g0635(.A(new_n829), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n631), .A2(new_n634), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n631), .A2(new_n634), .A3(new_n836), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT100), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n828), .B1(new_n740), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n684), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n627), .A2(new_n840), .A3(new_n682), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n727), .B1(new_n845), .B2(new_n709), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n709), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n841), .A2(new_n847), .ZN(G384));
  OAI21_X1  g0648(.A(new_n375), .B1(new_n360), .B2(new_n368), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT102), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n339), .A2(new_n648), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n358), .A2(KEYINPUT73), .A3(new_n359), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n366), .A2(new_n367), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT102), .B1(new_n857), .B2(new_n851), .ZN(new_n858));
  INV_X1    g0658(.A(new_n376), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n636), .A2(new_n852), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n853), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n707), .A2(new_n704), .A3(new_n705), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n861), .A2(new_n842), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n646), .B(KEYINPUT104), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n439), .B1(new_n438), .B2(new_n867), .ZN(new_n868));
  AND4_X1   g0668(.A1(new_n866), .A2(new_n868), .A3(new_n429), .A4(new_n430), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT16), .B1(new_n386), .B2(new_n391), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT103), .B1(new_n870), .B2(new_n287), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n380), .A3(new_n382), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n390), .B1(new_n874), .B2(G68), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n872), .B(new_n282), .C1(new_n875), .C2(KEYINPUT16), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n392), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n401), .ZN(new_n878));
  INV_X1    g0678(.A(new_n646), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n438), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n429), .A2(new_n430), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n869), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n432), .B2(new_n442), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n865), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n866), .A3(new_n868), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n646), .B1(new_n877), .B2(new_n401), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n437), .B1(new_n877), .B2(new_n401), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n429), .A2(new_n430), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n891), .B2(new_n866), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n443), .A2(new_n888), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(KEYINPUT38), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT105), .B(new_n865), .C1(new_n884), .C2(new_n885), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT106), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n864), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n867), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n422), .B(new_n903), .C1(new_n432), .C2(new_n442), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n427), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n422), .A2(KEYINPUT107), .A3(new_n413), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n868), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n869), .B1(KEYINPUT37), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n865), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n894), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n864), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n377), .A2(new_n443), .A3(new_n863), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n326), .A2(new_n648), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n844), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n861), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n898), .B2(new_n899), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n896), .A2(new_n897), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n376), .A2(new_n682), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n910), .B2(new_n894), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n903), .B1(new_n440), .B2(new_n441), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n922), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n444), .B1(new_n683), .B2(new_n685), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n641), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n931), .B(new_n933), .Z(new_n934));
  OAI22_X1  g0734(.A1(new_n917), .A2(new_n934), .B1(new_n245), .B2(new_n721), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n917), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n213), .A4(new_n448), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n387), .A2(new_n214), .A3(new_n260), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT101), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n941), .A2(new_n942), .B1(new_n202), .B2(G68), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n245), .B(G13), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n936), .A2(new_n940), .A3(new_n945), .ZN(G367));
  AOI211_X1 g0746(.A(new_n675), .B(new_n674), .C1(new_n573), .C2(new_n648), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n590), .A2(new_n682), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n949), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT42), .B1(new_n949), .B2(new_n661), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n532), .A3(new_n555), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n590), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n950), .A2(new_n951), .B1(new_n648), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT109), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n610), .A2(new_n682), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n680), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n612), .B2(new_n956), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT108), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT43), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n959), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n955), .B(new_n960), .C1(new_n962), .C2(new_n954), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n949), .A2(new_n654), .A3(new_n658), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n949), .A2(new_n662), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n659), .A2(KEYINPUT110), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n949), .A2(new_n662), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n659), .A2(KEYINPUT110), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n970), .B(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n967), .B(KEYINPUT45), .ZN(new_n976));
  OAI211_X1 g0776(.A(KEYINPUT110), .B(new_n659), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n658), .A2(new_n660), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n661), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n654), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n710), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n713), .B(KEYINPUT41), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n722), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n966), .A2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n743), .B1(new_n208), .B2(new_n316), .C1(new_n734), .C2(new_n233), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n727), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n766), .A2(new_n448), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n989), .A2(KEYINPUT46), .B1(new_n306), .B2(new_n778), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n378), .B1(new_n785), .B2(new_n822), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G294), .C2(new_n762), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n775), .A2(new_n462), .B1(new_n770), .B2(new_n815), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(KEYINPUT46), .B2(new_n989), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT111), .B(G317), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n994), .C1(new_n755), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G97), .B2(new_n752), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT112), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n752), .A2(G77), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n257), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n806), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G150), .A2(new_n774), .B1(new_n771), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n330), .B2(new_n778), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n766), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G50), .A2(new_n768), .B1(new_n1004), .B2(G58), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n790), .B2(new_n763), .C1(new_n805), .C2(new_n755), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1000), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n999), .A2(new_n998), .A3(new_n257), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n997), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  AOI21_X1  g0810(.A(new_n988), .B1(new_n1010), .B2(new_n742), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n962), .A2(new_n741), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n986), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n982), .A2(new_n723), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n658), .A2(new_n796), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n779), .A2(new_n500), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n775), .B2(new_n202), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n257), .B1(new_n770), .B2(new_n790), .C1(new_n785), .C2(new_n330), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n276), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1019), .C1(new_n1020), .C2(new_n762), .ZN(new_n1021));
  INV_X1    g0821(.A(G150), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n755), .A2(new_n1022), .B1(new_n260), .B2(new_n766), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT115), .Z(new_n1024));
  INV_X1    g0824(.A(new_n752), .ZN(new_n1025));
  INV_X1    g0825(.A(G97), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1021), .B(new_n1024), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G303), .A2(new_n768), .B1(new_n762), .B2(G311), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n776), .B2(new_n770), .C1(new_n775), .C2(new_n995), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1004), .A2(G294), .B1(new_n779), .B2(G283), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT117), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n755), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n257), .B1(new_n1038), .B2(G326), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(new_n448), .C2(new_n1025), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1036), .A2(KEYINPUT117), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1027), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n742), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n230), .A2(new_n250), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n271), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n717), .C1(G68), .C2(G77), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n734), .B(new_n1044), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n717), .A2(new_n208), .A3(new_n257), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(G107), .B2(new_n208), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n743), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1043), .A2(new_n727), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n982), .A2(new_n686), .A3(new_n709), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n713), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n982), .B1(new_n686), .B2(new_n709), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1015), .B1(new_n1016), .B2(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  INV_X1    g0858(.A(new_n1055), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n714), .B1(new_n978), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n973), .A2(new_n977), .A3(new_n1055), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n978), .A2(new_n723), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n775), .A2(new_n790), .B1(new_n770), .B2(new_n1022), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1038), .A2(new_n1001), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n257), .B1(new_n785), .B2(new_n271), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n763), .A2(new_n202), .B1(new_n330), .B2(new_n766), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G77), .C2(new_n779), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n817), .A2(new_n1065), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n378), .B1(new_n763), .B2(new_n462), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n785), .A2(new_n820), .B1(new_n766), .B2(new_n822), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G116), .C2(new_n779), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n782), .B(new_n1073), .C1(new_n776), .C2(new_n755), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n774), .B1(new_n771), .B2(G317), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1070), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n742), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n733), .A2(new_n237), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n744), .B1(G97), .B2(new_n712), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n726), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(new_n949), .C2(new_n796), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1063), .A2(KEYINPUT118), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT118), .B1(new_n1063), .B2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1062), .B1(new_n1083), .B2(new_n1084), .ZN(G390));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n668), .A2(new_n669), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n675), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n590), .A2(new_n596), .A3(new_n673), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n678), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n559), .B(new_n612), .C1(new_n625), .C2(KEYINPUT88), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n680), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n682), .B(new_n840), .C1(new_n1087), .C2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n862), .A2(G330), .A3(new_n840), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n861), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1095), .A3(new_n919), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n708), .A2(G330), .A3(new_n840), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n861), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n861), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n853), .A2(new_n858), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n859), .A2(new_n860), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n862), .A2(G330), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n840), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n920), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n444), .A2(new_n1104), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n932), .A2(new_n641), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1086), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n932), .A2(new_n641), .A3(new_n1108), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n861), .A2(new_n1094), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n861), .B2(new_n1097), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1113), .A2(new_n920), .B1(new_n1098), .B2(new_n1096), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT119), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1093), .A2(new_n919), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n925), .B(new_n911), .C1(new_n1118), .C2(new_n861), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n927), .B1(new_n923), .B2(KEYINPUT39), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n921), .A2(new_n926), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1112), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1119), .B1(new_n861), .B2(new_n1097), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1116), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n713), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n727), .B1(new_n1020), .B2(new_n801), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1120), .A2(new_n740), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n774), .A2(G116), .B1(G77), .B2(new_n779), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n822), .B2(new_n770), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n785), .A2(new_n1026), .B1(new_n763), .B2(new_n306), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n257), .A4(new_n788), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n811), .B(new_n1135), .C1(new_n820), .C2(new_n758), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT120), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n752), .A2(G50), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n759), .A2(G125), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1004), .A2(G150), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT53), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G128), .B2(new_n771), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n257), .B1(new_n763), .B2(new_n805), .ZN(new_n1144));
  INV_X1    g0944(.A(G132), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n775), .A2(new_n1145), .B1(new_n778), .B2(new_n790), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1144), .B(new_n1146), .C1(new_n768), .C2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1139), .A2(new_n1140), .A3(new_n1143), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1138), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1130), .B(new_n1131), .C1(new_n742), .C2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n723), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1129), .A2(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1128), .B2(new_n1111), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n290), .A2(new_n646), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n304), .B(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n912), .A2(G330), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n902), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1162), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1163), .B(new_n1166), .C1(new_n900), .C2(new_n901), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n931), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT106), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n923), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n896), .A2(KEYINPUT106), .A3(new_n897), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT40), .B1(new_n1173), .B2(new_n864), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1166), .B1(new_n1174), .B2(new_n1163), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n902), .A2(new_n1164), .A3(new_n1162), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n931), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1158), .B1(new_n1169), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n713), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT122), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n931), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n922), .A2(new_n929), .A3(KEYINPUT122), .A4(new_n930), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1175), .A2(new_n1176), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1168), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1128), .A2(new_n1111), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1179), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n752), .A2(G58), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n257), .B(new_n471), .C1(new_n1004), .C2(G77), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(new_n822), .C2(new_n758), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT121), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n775), .A2(new_n306), .B1(new_n770), .B2(new_n448), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1026), .A2(new_n763), .B1(new_n785), .B2(new_n316), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G68), .C2(new_n779), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(KEYINPUT58), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G33), .A2(G41), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G50), .B(new_n1197), .C1(new_n378), .C2(new_n342), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1038), .A2(G124), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n1025), .C2(new_n790), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n774), .A2(G128), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1022), .B2(new_n778), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G125), .B2(new_n771), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G132), .A2(new_n762), .B1(new_n1004), .B2(new_n1148), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n805), .C2(new_n785), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1200), .B1(KEYINPUT59), .B2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1198), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1196), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT58), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n742), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n727), .C1(G50), .C2(new_n801), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n739), .B2(new_n1162), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1185), .B2(new_n723), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1188), .A2(new_n1214), .ZN(G375));
  OAI22_X1  g1015(.A1(new_n1147), .A2(new_n763), .B1(new_n785), .B2(new_n1022), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n378), .B(new_n1216), .C1(G159), .C2(new_n1004), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n759), .A2(G128), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n770), .A2(new_n1145), .B1(new_n778), .B2(new_n202), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G137), .B2(new_n774), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1189), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n763), .A2(new_n448), .B1(new_n1026), .B2(new_n766), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n257), .B(new_n1222), .C1(G107), .C2(new_n768), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1017), .B1(new_n820), .B2(new_n770), .C1(new_n775), .C2(new_n822), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n999), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n758), .A2(new_n462), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n742), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n726), .B1(new_n330), .B2(new_n800), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n1103), .C2(new_n740), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1107), .B2(new_n722), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT123), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n984), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1116), .B2(new_n1236), .ZN(G381));
  OR3_X1    g1037(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1239), .A2(new_n1188), .A3(new_n1240), .A4(new_n1214), .ZN(G407));
  NAND2_X1  g1041(.A1(new_n647), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G375), .C2(new_n1244), .ZN(G409));
  INV_X1    g1045(.A(KEYINPUT127), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n966), .A2(new_n985), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G390), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(G390), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1247), .B2(G390), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(G393), .B(new_n798), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n1249), .A2(new_n1250), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1247), .A2(G390), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1256), .A2(new_n1251), .A3(new_n1248), .A4(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1214), .C1(new_n1179), .C2(new_n1187), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1175), .A2(new_n931), .A3(new_n1176), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1184), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1213), .B1(new_n1263), .B2(new_n723), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1185), .A2(new_n1235), .A3(new_n1186), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1240), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1243), .B1(new_n1261), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n713), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1110), .A2(new_n1115), .A3(KEYINPUT60), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1234), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(G384), .A3(new_n1233), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  XOR2_X1   g1075(.A(new_n1232), .B(KEYINPUT123), .Z(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1272), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1243), .A2(G2897), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1284), .B2(new_n1280), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1260), .B1(new_n1268), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G384), .B1(new_n1273), .B2(new_n1233), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1276), .A2(new_n1272), .A3(new_n1275), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1268), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1286), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1268), .A2(new_n1287), .A3(new_n1290), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1259), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1261), .A2(new_n1267), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1242), .A3(new_n1290), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1255), .A2(new_n1260), .A3(new_n1257), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT125), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1280), .B1(new_n1302), .B2(new_n1279), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1281), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1268), .B2(KEYINPUT124), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1295), .A2(KEYINPUT124), .A3(new_n1242), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1301), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1246), .B1(new_n1294), .B2(new_n1309), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1268), .A2(new_n1285), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1260), .A4(new_n1293), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1258), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1255), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1297), .B2(new_n1296), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1316), .B(new_n1299), .C1(new_n1307), .C2(new_n1306), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1317), .A3(KEYINPUT127), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1240), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1261), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1290), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1258), .ZN(G402));
endmodule


