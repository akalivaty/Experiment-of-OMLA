//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n203), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n201), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n222), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G58), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n213), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n213), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n213), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n249), .B1(new_n250), .B2(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n212), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n255), .A2(new_n260), .B1(new_n246), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n257), .A2(new_n259), .A3(new_n212), .A4(new_n262), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G226), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n270), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT65), .B(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n277), .B(new_n261), .C1(new_n278), .C2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G222), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G223), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n283), .B1(new_n284), .B2(new_n281), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n280), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n269), .B(new_n291), .C1(G169), .C2(new_n289), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n268), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT68), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n269), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n294), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n294), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n305), .A2(new_n307), .A3(G226), .A4(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G87), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n307), .A3(G223), .A4(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n281), .A2(KEYINPUT73), .A3(G223), .A4(new_n282), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n304), .B1(new_n315), .B2(new_n271), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n279), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n313), .A2(new_n314), .ZN(new_n323));
  INV_X1    g0123(.A(new_n310), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n318), .B1(new_n325), .B2(new_n288), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n316), .A2(new_n322), .B1(new_n326), .B2(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n305), .A2(new_n307), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n328), .B2(new_n213), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT7), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n330), .B(G20), .C1(new_n305), .C2(new_n307), .ZN(new_n331));
  OAI21_X1  g0131(.A(G68), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n334), .B2(new_n245), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G20), .A2(G33), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G159), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n213), .B1(new_n203), .B2(new_n333), .ZN(new_n340));
  INV_X1    g0140(.A(new_n338), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT71), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n330), .B1(new_n281), .B2(G20), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n202), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n335), .A2(new_n338), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n343), .A2(new_n349), .A3(new_n260), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n254), .A2(new_n263), .ZN(new_n351));
  XOR2_X1   g0151(.A(KEYINPUT8), .B(G58), .Z(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n267), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(new_n265), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT72), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n354), .B(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n327), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT17), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n350), .A2(new_n356), .ZN(new_n360));
  INV_X1    g0160(.A(new_n321), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT74), .B1(new_n279), .B2(new_n317), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(G179), .B1(new_n325), .B2(new_n288), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n279), .A2(new_n317), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n315), .B2(new_n271), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n363), .A2(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT18), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n327), .A2(KEYINPUT17), .A3(new_n350), .A4(new_n356), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n359), .A2(new_n370), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n273), .A2(G238), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n376), .A2(new_n279), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n281), .A2(G232), .A3(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G97), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n305), .A2(new_n307), .A3(G226), .A4(new_n282), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n288), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n377), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g0185(.A(G169), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n382), .A2(new_n288), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n376), .A2(new_n279), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT69), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT69), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT13), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n377), .A2(new_n383), .A3(new_n378), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(G169), .C1(new_n384), .C2(new_n385), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n387), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n253), .A2(new_n284), .B1(new_n213), .B2(G68), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n400), .A2(KEYINPUT70), .B1(new_n246), .B2(new_n252), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n260), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT11), .B(new_n260), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n263), .A2(new_n202), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT12), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n266), .A2(G68), .A3(new_n267), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n393), .A2(G190), .A3(new_n394), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT13), .B1(new_n388), .B2(new_n389), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n394), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(G200), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n399), .A2(new_n410), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n352), .A2(new_n337), .B1(G20), .B2(G77), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n253), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n260), .B1(new_n284), .B2(new_n263), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n266), .A2(G77), .A3(new_n267), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n281), .A2(G232), .A3(new_n282), .ZN(new_n422));
  INV_X1    g0222(.A(G107), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n423), .B2(new_n281), .C1(new_n285), .C2(new_n217), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n288), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n273), .A2(G244), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n279), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n421), .B1(new_n429), .B2(G190), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n297), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n290), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n428), .A2(new_n367), .B1(new_n419), .B2(new_n420), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n375), .A2(new_n415), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n303), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G45), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n219), .B1(new_n438), .B2(G1), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n261), .A2(new_n275), .A3(G45), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n271), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(G1698), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n305), .A2(new_n307), .A3(G238), .A4(new_n282), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G116), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI211_X1 g0245(.A(G179), .B(new_n441), .C1(new_n445), .C2(new_n288), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n288), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n367), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n265), .B1(new_n261), .B2(G33), .ZN(new_n450));
  INV_X1    g0250(.A(new_n417), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT19), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n213), .B1(new_n380), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G97), .A2(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n218), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n305), .A2(new_n307), .A3(new_n213), .A4(G68), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n253), .B2(new_n223), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n260), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n417), .A2(new_n263), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n304), .B(new_n441), .C1(new_n445), .C2(new_n288), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n257), .A2(new_n212), .A3(new_n259), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n261), .A2(G33), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(G87), .A3(new_n262), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n467), .A3(new_n462), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n448), .A2(G200), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n449), .A2(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n329), .B2(new_n331), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n423), .A2(KEYINPUT6), .A3(G97), .ZN(new_n473));
  AND2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n455), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(KEYINPUT6), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(G20), .B1(G77), .B2(new_n337), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n260), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n450), .A2(G97), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n262), .A2(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(new_n282), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G283), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n251), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G250), .A2(G1698), .ZN(new_n489));
  NAND2_X1  g0289(.A1(KEYINPUT4), .A2(G244), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G1698), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n281), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n271), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT75), .B1(new_n495), .B2(G41), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT75), .ZN(new_n497));
  INV_X1    g0297(.A(G41), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT5), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT65), .A2(G41), .ZN(new_n501));
  NOR2_X1   g0301(.A1(KEYINPUT65), .A2(G41), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n438), .A2(G1), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n500), .A2(new_n277), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(G257), .A3(new_n271), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n494), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n367), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n507), .A2(G257), .A3(new_n271), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n277), .A2(new_n499), .A3(new_n496), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n503), .A2(new_n504), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n511), .A2(new_n493), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n290), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n483), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n494), .A2(new_n304), .A3(new_n505), .A4(new_n508), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n515), .B2(G200), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n465), .B1(new_n472), .B2(new_n477), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n450), .A2(G97), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(new_n481), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n471), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n266), .A2(G116), .A3(new_n466), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n263), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n251), .A2(G97), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(G20), .B2(new_n526), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n260), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n525), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n271), .B1(new_n328), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(G257), .A2(G1698), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n282), .A2(G264), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n281), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n535), .A2(KEYINPUT76), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT76), .B1(new_n535), .B2(new_n538), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n507), .A2(G270), .A3(new_n271), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n505), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n541), .A2(new_n543), .A3(new_n290), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT21), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n367), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n542), .A2(new_n505), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT76), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n537), .A2(new_n536), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n328), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n288), .B1(new_n281), .B2(G303), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n535), .A2(KEYINPUT76), .A3(new_n538), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n547), .B1(new_n548), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n533), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n533), .B(G169), .C1(new_n541), .C2(new_n543), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  INV_X1    g0359(.A(new_n533), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n548), .A2(G190), .A3(new_n555), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n541), .A2(new_n543), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(new_n297), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n557), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT80), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n305), .A2(new_n307), .A3(new_n213), .A4(G87), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n281), .A2(KEYINPUT22), .A3(new_n213), .A4(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT77), .B1(new_n444), .B2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT77), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n573), .A2(new_n213), .A3(G33), .A4(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT78), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n213), .C2(G107), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n213), .A2(G107), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT79), .B1(new_n581), .B2(new_n577), .ZN(new_n582));
  AND4_X1   g0382(.A1(KEYINPUT79), .A2(new_n577), .A3(new_n423), .A4(G20), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n575), .B(new_n580), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n565), .B(new_n566), .C1(new_n571), .C2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n565), .B1(new_n571), .B2(new_n584), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n576), .A2(new_n577), .B1(new_n423), .B2(G20), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n579), .A2(new_n590), .B1(new_n572), .B2(new_n574), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n569), .A4(new_n570), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n565), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n260), .B(new_n585), .C1(new_n587), .C2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n266), .A2(G107), .A3(new_n466), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n263), .A2(new_n423), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT25), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT81), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n450), .A2(G107), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT25), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n596), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n507), .A2(G264), .A3(new_n271), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n219), .A2(new_n282), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n224), .A2(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n305), .A2(new_n606), .A3(new_n307), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n288), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n611), .A3(new_n505), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT82), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n605), .A2(new_n611), .A3(new_n614), .A4(new_n505), .ZN(new_n615));
  AOI21_X1  g0415(.A(G190), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n612), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n594), .B(new_n604), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(G169), .A3(new_n615), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(G179), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n585), .A2(new_n260), .ZN(new_n623));
  INV_X1    g0423(.A(new_n593), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n566), .B1(new_n592), .B2(new_n565), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n604), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n524), .A2(new_n564), .A3(new_n619), .A4(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n437), .A2(new_n629), .ZN(G372));
  NAND2_X1  g0430(.A1(new_n399), .A2(new_n410), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n414), .A2(new_n411), .ZN(new_n632));
  INV_X1    g0432(.A(new_n434), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n635), .A2(new_n359), .A3(new_n373), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n370), .A2(new_n372), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n636), .A2(new_n638), .B1(new_n302), .B2(new_n301), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n292), .ZN(new_n640));
  INV_X1    g0440(.A(new_n517), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .A3(new_n471), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n449), .A2(new_n463), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n469), .A2(new_n470), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n517), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n644), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n594), .A2(new_n604), .B1(new_n620), .B2(new_n621), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n557), .A2(new_n559), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n524), .B(new_n619), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n640), .B1(new_n437), .B2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n557), .A2(new_n563), .A3(new_n559), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT83), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n261), .A2(new_n213), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n560), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n656), .B2(KEYINPUT83), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n546), .B1(new_n541), .B2(new_n543), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n548), .A2(G179), .A3(new_n555), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n669), .A2(new_n533), .B1(new_n558), .B2(new_n545), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n657), .A2(new_n666), .B1(new_n670), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n628), .A2(new_n619), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n664), .B1(new_n594), .B2(new_n604), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n628), .B2(new_n664), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n663), .B(KEYINPUT84), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n650), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n674), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n651), .A2(new_n664), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n677), .A2(new_n679), .A3(new_n683), .ZN(G399));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n605), .A2(new_n611), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT85), .B1(new_n448), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT85), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n447), .A2(new_n688), .A3(new_n605), .A4(new_n611), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n544), .A2(new_n687), .A3(new_n515), .A4(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n562), .A2(new_n515), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n290), .A3(new_n612), .A4(new_n448), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n509), .A2(new_n691), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n544), .A3(new_n687), .A4(new_n689), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n692), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n678), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT86), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n697), .A2(KEYINPUT86), .A3(KEYINPUT31), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n663), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT87), .B1(new_n629), .B2(new_n698), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n471), .A2(new_n517), .A3(new_n523), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n656), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT87), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n680), .A2(new_n709), .A3(new_n710), .A4(new_n678), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n685), .B1(new_n706), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT88), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI211_X1 g0515(.A(KEYINPUT88), .B(new_n685), .C1(new_n706), .C2(new_n712), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n698), .B1(new_n649), .B2(new_n652), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n653), .B2(new_n664), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(KEYINPUT89), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n711), .B2(new_n707), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT88), .B1(new_n725), .B2(new_n685), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n713), .A2(new_n714), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT89), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n723), .A2(new_n730), .A3(new_n261), .ZN(new_n731));
  INV_X1    g0531(.A(new_n207), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n278), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n456), .A2(G116), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n210), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(new_n738), .ZN(G364));
  INV_X1    g0539(.A(G13), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n261), .B1(new_n741), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n673), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n671), .A2(G330), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT90), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n671), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n281), .A2(new_n207), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n207), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n240), .A2(new_n438), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n732), .A2(new_n281), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n438), .B2(new_n211), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n755), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n212), .B1(G20), .B2(new_n367), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n744), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n213), .B1(new_n765), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(G294), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n213), .A2(G190), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n290), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n328), .B1(new_n766), .B2(new_n767), .C1(new_n768), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n213), .A2(new_n304), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n770), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n765), .ZN(new_n776));
  INV_X1    g0576(.A(G329), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n290), .A2(new_n297), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n769), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n779), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n772), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n769), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(G179), .A3(new_n297), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT91), .Z(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n773), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(new_n297), .A3(G179), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT93), .Z(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n785), .B1(new_n789), .B2(new_n487), .C1(new_n534), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n788), .A2(G107), .ZN(new_n795));
  INV_X1    g0595(.A(new_n791), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n281), .C1(new_n218), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT92), .ZN(new_n798));
  INV_X1    g0598(.A(new_n780), .ZN(new_n799));
  INV_X1    g0599(.A(new_n771), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G68), .A2(new_n799), .B1(new_n800), .B2(G77), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n801), .B1(new_n246), .B2(new_n782), .C1(new_n201), .C2(new_n774), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n766), .A2(new_n223), .ZN(new_n803));
  INV_X1    g0603(.A(new_n776), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G159), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  OR3_X1    g0606(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n794), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n764), .B1(new_n808), .B2(new_n761), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n745), .A2(new_n747), .B1(new_n752), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NOR2_X1   g0611(.A1(new_n434), .A2(new_n663), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n421), .A2(new_n663), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n431), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n434), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n718), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n717), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT95), .Z(new_n818));
  AOI21_X1  g0618(.A(new_n744), .B1(new_n717), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n744), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n761), .A2(new_n748), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n284), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n281), .B1(new_n766), .B2(new_n201), .C1(new_n824), .C2(new_n776), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n789), .A2(new_n202), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G50), .C2(new_n792), .ZN(new_n827));
  INV_X1    g0627(.A(new_n774), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G143), .A2(new_n828), .B1(new_n800), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n782), .C1(new_n250), .C2(new_n780), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT34), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n782), .A2(new_n534), .B1(new_n780), .B2(new_n487), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G116), .B2(new_n800), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT94), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n788), .A2(G87), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n793), .B2(new_n423), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n328), .B1(new_n776), .B2(new_n768), .C1(new_n767), .C2(new_n774), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n837), .A2(new_n803), .A3(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n827), .A2(new_n832), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n761), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n823), .B1(new_n840), .B2(new_n841), .C1(new_n815), .C2(new_n749), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n820), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n741), .A2(new_n261), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT40), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  INV_X1    g0646(.A(new_n661), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n360), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n357), .A2(new_n369), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n342), .A2(new_n339), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n347), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n465), .B1(new_n853), .B2(KEYINPUT16), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n344), .B1(new_n852), .B2(new_n347), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n354), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n290), .B1(new_n315), .B2(new_n271), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n322), .A2(new_n857), .B1(new_n326), .B2(G169), .ZN(new_n858));
  AOI21_X1  g0658(.A(G190), .B1(new_n325), .B2(new_n288), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n363), .A2(new_n859), .B1(new_n366), .B2(new_n297), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n856), .A2(new_n858), .B1(new_n360), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT97), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT97), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n357), .B(new_n863), .C1(new_n858), .C2(new_n856), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n856), .A2(new_n661), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n851), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n374), .A2(new_n865), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n846), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n865), .B1(new_n861), .B2(KEYINPUT97), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n849), .B1(new_n872), .B2(new_n864), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n869), .B(KEYINPUT38), .C1(new_n873), .C2(new_n851), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n410), .A2(new_n663), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI221_X4 g0677(.A(new_n877), .B1(new_n411), .B2(new_n414), .C1(new_n399), .C2(new_n410), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n631), .B2(new_n632), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n815), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT31), .B1(new_n697), .B2(new_n663), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n712), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n875), .B1(new_n884), .B2(KEYINPUT99), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n674), .A2(new_n708), .A3(new_n656), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n710), .B1(new_n886), .B2(new_n678), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n481), .B1(new_n478), .B2(new_n260), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n480), .B1(new_n290), .B2(new_n515), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n510), .B1(new_n522), .B2(new_n519), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n890), .A2(new_n471), .A3(new_n670), .A4(new_n563), .ZN(new_n891));
  NOR4_X1   g0691(.A1(new_n891), .A2(new_n674), .A3(KEYINPUT87), .A4(new_n698), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n883), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n880), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n845), .B1(new_n885), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n357), .A2(new_n369), .A3(new_n848), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n850), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT98), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT98), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n901), .A3(new_n850), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n374), .A2(new_n360), .A3(new_n847), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n846), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n845), .B1(new_n905), .B2(new_n874), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n884), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n436), .A2(new_n893), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT101), .Z(new_n911));
  AOI21_X1  g0711(.A(new_n685), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n878), .A2(new_n879), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n648), .A2(new_n644), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n628), .A2(new_n670), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n917), .A2(new_n524), .A3(new_n619), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n678), .B(new_n815), .C1(new_n916), .C2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n812), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n875), .A2(new_n915), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n638), .A2(new_n661), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT39), .B1(new_n905), .B2(new_n874), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n631), .A2(new_n663), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n436), .B1(new_n720), .B2(new_n721), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n640), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n931), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n844), .B1(new_n913), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n913), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n476), .B(KEYINPUT96), .Z(new_n937));
  INV_X1    g0737(.A(KEYINPUT35), .ZN(new_n938));
  OAI211_X1 g0738(.A(G116), .B(new_n214), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n937), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT36), .Z(new_n941));
  NAND3_X1  g0741(.A1(new_n211), .A2(G77), .A3(new_n333), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(G50), .B2(new_n202), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n740), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT102), .Z(G367));
  OR2_X1    g0746(.A1(new_n236), .A2(new_n758), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n763), .B1(new_n732), .B2(new_n451), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n821), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n468), .A2(new_n663), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n644), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n471), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n787), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n954), .A2(new_n284), .B1(new_n776), .B2(new_n830), .ZN(new_n955));
  INV_X1    g0755(.A(G159), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n780), .A2(new_n956), .B1(new_n771), .B2(new_n246), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT107), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n796), .A2(new_n201), .B1(new_n774), .B2(new_n250), .ZN(new_n959));
  INV_X1    g0759(.A(G143), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n281), .B1(new_n766), .B2(new_n202), .C1(new_n782), .C2(new_n960), .ZN(new_n961));
  OR4_X1    g0761(.A1(new_n955), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT105), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n767), .A2(new_n780), .B1(new_n774), .B2(new_n534), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT46), .B1(new_n791), .B2(G116), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT106), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n782), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n965), .B(new_n968), .C1(G311), .C2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n328), .B1(new_n771), .B2(new_n487), .ZN(new_n971));
  INV_X1    g0771(.A(G317), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n954), .A2(new_n223), .B1(new_n776), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n766), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n971), .B(new_n973), .C1(G107), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n966), .A2(new_n967), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n962), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI221_X1 g0779(.A(new_n949), .B1(new_n751), .B2(new_n953), .C1(new_n979), .C2(new_n841), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n683), .A2(new_n679), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n641), .A2(new_n698), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n517), .B(new_n523), .C1(new_n522), .C2(new_n678), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n982), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT44), .B1(new_n982), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n683), .A2(new_n679), .A3(new_n985), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT104), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n677), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n676), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n990), .A2(new_n993), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n994), .B(new_n677), .C1(new_n989), .C2(new_n992), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n672), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n723), .A2(new_n730), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n733), .B(KEYINPUT41), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n742), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n683), .A2(new_n986), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT103), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n517), .B1(new_n984), .B2(new_n628), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1008), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1006), .B(KEYINPUT103), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT42), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n953), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n677), .A2(new_n986), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1010), .A2(new_n1016), .A3(new_n1015), .A4(new_n1013), .ZN(new_n1021));
  AND3_X1   g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n981), .B1(new_n1005), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(G387));
  AOI21_X1  g0826(.A(KEYINPUT89), .B1(new_n717), .B2(new_n722), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n728), .A2(new_n729), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1002), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n723), .A2(new_n730), .A3(new_n1001), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1029), .A2(new_n733), .A3(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n676), .A2(new_n751), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n753), .A2(new_n735), .B1(G107), .B2(new_n207), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT108), .Z(new_n1034));
  OR2_X1    g0834(.A1(new_n232), .A2(new_n438), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n735), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n1036), .C1(G68), .C2(G77), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n254), .A2(G50), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n758), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n744), .B1(new_n1041), .B2(new_n763), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n788), .A2(G97), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n780), .A2(new_n254), .B1(new_n771), .B2(new_n202), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n774), .A2(new_n246), .B1(new_n776), .B2(new_n250), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n796), .A2(new_n284), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n766), .A2(new_n417), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n328), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n969), .A2(G159), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT109), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1043), .A2(new_n1046), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n796), .A2(new_n767), .B1(new_n766), .B2(new_n487), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n828), .B1(new_n800), .B2(G303), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n768), .B2(new_n780), .C1(new_n775), .C2(new_n782), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT49), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n328), .B1(new_n783), .B2(new_n776), .C1(new_n954), .C2(new_n526), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1042), .B1(new_n1061), .B2(new_n761), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1002), .A2(new_n743), .B1(new_n1032), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1031), .A2(new_n1063), .ZN(G393));
  NAND2_X1  g0864(.A1(new_n999), .A2(new_n743), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n762), .B1(new_n223), .B2(new_n207), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n243), .A2(new_n758), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n744), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n796), .A2(new_n487), .B1(new_n780), .B2(new_n534), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G294), .B2(new_n800), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n328), .B1(new_n776), .B2(new_n775), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G116), .B2(new_n974), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n795), .A3(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n782), .A2(new_n972), .B1(new_n774), .B2(new_n768), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n782), .A2(new_n250), .B1(new_n774), .B2(new_n956), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n281), .B1(new_n776), .B2(new_n960), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n791), .B2(G68), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n836), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n780), .A2(new_n246), .B1(new_n771), .B2(new_n254), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n766), .A2(new_n284), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT110), .Z(new_n1084));
  OAI22_X1  g0884(.A1(new_n1073), .A2(new_n1075), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1068), .B1(new_n1085), .B2(new_n761), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n985), .B2(new_n751), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1065), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1001), .B1(new_n723), .B2(new_n730), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n999), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n733), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1090), .A2(new_n999), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n726), .A2(new_n727), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n815), .A3(new_n915), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n921), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n914), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n929), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1098), .A2(new_n928), .B1(new_n1099), .B2(new_n926), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n814), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n633), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n663), .B(new_n1102), .C1(new_n649), .C2(new_n652), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n915), .B1(new_n1103), .B2(new_n812), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n905), .A2(new_n874), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n928), .B(KEYINPUT111), .Z(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1096), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n893), .A2(G330), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(new_n880), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n928), .B1(new_n921), .B2(new_n915), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n927), .B2(new_n929), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n932), .B(new_n640), .C1(new_n437), .C2(new_n1109), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n893), .A2(G330), .A3(new_n815), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n812), .B(new_n1103), .C1(new_n1118), .C2(new_n914), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n815), .B1(new_n715), .B2(new_n716), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1110), .B1(new_n1121), .B2(new_n914), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n1097), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1115), .A2(new_n1117), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n815), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n726), .B2(new_n727), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(new_n915), .B1(new_n880), .B2(new_n1109), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1128), .A2(new_n921), .B1(new_n1096), .B2(new_n1119), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1125), .B1(new_n1129), .B2(new_n1116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1124), .A2(new_n1130), .A3(new_n733), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n826), .B1(G87), .B2(new_n792), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G116), .A2(new_n828), .B1(new_n800), .B2(G97), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n969), .A2(G283), .B1(new_n804), .B2(G294), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n281), .B(new_n1082), .C1(G107), .C2(new_n799), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n791), .A2(G150), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT113), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT53), .Z(new_n1139));
  AOI22_X1  g0939(.A1(G128), .A2(new_n969), .B1(new_n828), .B2(G132), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT112), .Z(new_n1141));
  NOR2_X1   g0941(.A1(new_n954), .A2(new_n246), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n780), .A2(new_n830), .B1(new_n776), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT54), .B(G143), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n281), .B1(new_n766), .B2(new_n956), .C1(new_n771), .C2(new_n1145), .ZN(new_n1146));
  OR4_X1    g0946(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1136), .B1(new_n1139), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n761), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n822), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n744), .C1(new_n352), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n927), .A2(new_n929), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n749), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT114), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n743), .B2(new_n1115), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1131), .A2(new_n1156), .ZN(G378));
  NAND3_X1  g0957(.A1(new_n303), .A2(new_n269), .A3(new_n847), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n269), .A2(new_n847), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n292), .B(new_n1159), .C1(new_n301), .C2(new_n302), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(new_n749), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n223), .A2(new_n780), .B1(new_n774), .B2(new_n423), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1047), .A2(new_n281), .A3(new_n278), .A4(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n782), .A2(new_n526), .B1(new_n766), .B2(new_n202), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT115), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n804), .A2(G283), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n954), .A2(new_n201), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n451), .B2(new_n800), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n782), .A2(new_n1143), .B1(new_n780), .B2(new_n824), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1145), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n791), .A2(new_n1177), .B1(G128), .B2(new_n828), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n250), .B2(new_n766), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G137), .C2(new_n800), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n251), .B(new_n498), .C1(new_n954), .C2(new_n956), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G124), .B2(new_n804), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n246), .B1(G33), .B2(G41), .C1(new_n281), .C2(new_n278), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1188));
  AND4_X1   g0988(.A1(new_n1175), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n744), .B1(G50), .B2(new_n1150), .C1(new_n1189), .C2(new_n841), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1165), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1099), .A2(new_n926), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n924), .B1(new_n1192), .B2(new_n928), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n685), .B1(new_n906), .B2(new_n884), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n896), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n896), .B2(new_n1194), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT117), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n893), .A2(new_n894), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT99), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1201), .A2(new_n1202), .B1(new_n874), .B2(new_n871), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n884), .A2(KEYINPUT99), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT40), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n907), .A2(G330), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1164), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT116), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n896), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n925), .A2(new_n930), .A3(KEYINPUT117), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1200), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1191), .B1(new_n1215), .B2(new_n743), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1117), .B1(new_n1129), .B2(new_n1125), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1116), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1196), .A2(new_n1197), .A3(new_n1193), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n931), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1221));
  OAI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n733), .B1(new_n1219), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1216), .B1(new_n1218), .B2(new_n1223), .ZN(G375));
  OAI21_X1  g1024(.A(KEYINPUT118), .B1(new_n1129), .B2(new_n742), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT118), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1123), .A2(new_n1226), .A3(new_n743), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n914), .A2(new_n748), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n744), .B1(G68), .B2(new_n1150), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n780), .A2(new_n526), .B1(new_n771), .B2(new_n423), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n792), .A2(G97), .B1(KEYINPUT119), .B2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(KEYINPUT119), .B2(new_n1230), .C1(new_n284), .C2(new_n789), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n774), .A2(new_n487), .B1(new_n776), .B2(new_n534), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n328), .B1(new_n782), .B2(new_n767), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1048), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G132), .A2(new_n969), .B1(new_n799), .B2(new_n1177), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n830), .B2(new_n774), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT120), .Z(new_n1238));
  AOI211_X1 g1038(.A(new_n328), .B(new_n1171), .C1(G128), .C2(new_n804), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G150), .A2(new_n800), .B1(new_n974), .B2(G50), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT121), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT121), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n792), .A2(G159), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1232), .A2(new_n1235), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1229), .B1(new_n1245), .B2(new_n761), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT122), .Z(new_n1247));
  AOI22_X1  g1047(.A1(new_n1225), .A2(new_n1227), .B1(new_n1228), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1129), .A2(new_n1116), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1123), .A2(new_n1117), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1004), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(G381));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1029), .A2(new_n998), .A3(new_n997), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n734), .B1(new_n1090), .B2(new_n999), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1088), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1031), .A2(new_n810), .A3(new_n1063), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1025), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G378), .A2(G375), .A3(new_n1259), .A4(G381), .ZN(G407));
  XOR2_X1   g1060(.A(new_n1154), .B(KEYINPUT114), .Z(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n742), .B2(new_n1125), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n734), .B1(new_n1250), .B2(new_n1125), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1124), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n662), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G407), .B(G213), .C1(G375), .C2(new_n1267), .ZN(G409));
  XNOR2_X1  g1068(.A(new_n1025), .B(new_n1257), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(G390), .B2(new_n1025), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n810), .B1(new_n1031), .B2(new_n1063), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT125), .B1(new_n1258), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1031), .A2(new_n810), .A3(new_n1063), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1269), .A2(new_n1271), .A3(new_n1273), .A4(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1271), .A2(new_n1273), .A3(new_n1277), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G390), .B(new_n1025), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1214), .B1(new_n1221), .B2(KEYINPUT117), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1211), .B1(new_n1284), .B2(new_n1208), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1251), .B(new_n1217), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n743), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1191), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(KEYINPUT123), .A3(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT123), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1207), .A2(new_n931), .A3(new_n1209), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n742), .B1(new_n1198), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1292), .B2(new_n1191), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1286), .A2(new_n1289), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1264), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G378), .B(new_n1216), .C1(new_n1218), .C2(new_n1223), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1294), .B2(new_n1264), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1265), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n915), .B1(new_n1095), .B2(new_n815), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n921), .B1(new_n1301), .B2(new_n1110), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1302), .A2(KEYINPUT60), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n733), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1250), .A2(KEYINPUT60), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1249), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1247), .A2(new_n1228), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1129), .A2(KEYINPUT118), .A3(new_n742), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1226), .B1(new_n1123), .B2(new_n743), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1254), .B1(new_n1306), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1123), .B2(new_n1117), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1116), .B2(new_n1129), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1248), .B(G384), .C1(new_n1314), .C2(new_n1304), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1266), .A2(G2897), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1311), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1311), .B2(new_n1315), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI211_X1 g1119(.A(KEYINPUT61), .B(new_n1282), .C1(new_n1300), .C2(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1311), .A2(new_n1315), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1265), .B(new_n1321), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1299), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1266), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1327), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1321), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1320), .A2(new_n1324), .A3(new_n1328), .A4(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1319), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1326), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1333), .A2(new_n1334), .A3(new_n1265), .A4(new_n1321), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1322), .A2(KEYINPUT62), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1332), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1282), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1331), .A2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1264), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1282), .A2(new_n1340), .A3(new_n1297), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1297), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(new_n1278), .A3(new_n1281), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  XOR2_X1   g1144(.A(new_n1344), .B(new_n1321), .Z(G402));
endmodule


