//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n869, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G22gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G15gat), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G22gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(new_n205), .B2(new_n207), .ZN(new_n211));
  OAI21_X1  g010(.A(G8gat), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n208), .B(new_n213), .C1(new_n210), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G43gat), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(G43gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n218), .A2(G43gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n220), .A2(G50gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n229), .A2(new_n230), .A3(new_n224), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  OR3_X1    g032(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(G29gat), .B2(G36gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n231), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT17), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n236), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n231), .B1(new_n225), .B2(KEYINPUT87), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n228), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n243), .A2(new_n244), .A3(new_n238), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n216), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n212), .A2(new_n215), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n223), .A2(new_n227), .A3(new_n224), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n227), .B1(new_n223), .B2(new_n224), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n248), .A2(new_n249), .A3(new_n231), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n239), .B(new_n247), .C1(new_n250), .C2(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT89), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n238), .B1(new_n233), .B2(new_n236), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT88), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n246), .A2(new_n256), .A3(KEYINPUT18), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n253), .B2(new_n247), .ZN(new_n262));
  OAI211_X1 g061(.A(KEYINPUT91), .B(new_n216), .C1(new_n243), .C2(new_n238), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n252), .A2(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n258), .B(KEYINPUT13), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n239), .B1(new_n250), .B2(new_n241), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT91), .B1(new_n269), .B2(new_n216), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n253), .A2(new_n261), .A3(new_n247), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n254), .B1(new_n253), .B2(new_n247), .ZN(new_n272));
  NOR4_X1   g071(.A1(new_n243), .A2(KEYINPUT89), .A3(new_n238), .A4(new_n216), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT92), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  OAI211_X1 g074(.A(KEYINPUT90), .B(new_n260), .C1(new_n268), .C2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n246), .A2(new_n256), .A3(new_n259), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT18), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n260), .B(new_n279), .C1(new_n268), .C2(new_n275), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G141gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT11), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G197gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n285), .B(KEYINPUT12), .Z(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  AND4_X1   g086(.A1(KEYINPUT18), .A2(new_n246), .A3(new_n256), .A4(new_n259), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n265), .B1(new_n264), .B2(new_n267), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT92), .A3(new_n266), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n286), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n291), .B(new_n279), .C1(KEYINPUT90), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n296), .A2(KEYINPUT1), .ZN(new_n297));
  XOR2_X1   g096(.A(G127gat), .B(G134gat), .Z(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT71), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT72), .A4(new_n303), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G141gat), .B(G148gat), .Z(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT2), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G155gat), .B(G162gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT76), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n309), .A2(new_n317), .A3(new_n314), .A4(new_n312), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n316), .A2(new_n318), .B1(new_n315), .B2(new_n313), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n308), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n313), .A2(new_n315), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n307), .ZN(new_n327));
  INV_X1    g126(.A(new_n299), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n333));
  OAI211_X1 g132(.A(new_n322), .B(new_n332), .C1(new_n320), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n335), .ZN(new_n339));
  INV_X1    g138(.A(new_n320), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n308), .A2(new_n319), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT79), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(KEYINPUT5), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(new_n335), .ZN(new_n347));
  INV_X1    g146(.A(new_n333), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT78), .B1(new_n320), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n320), .A2(KEYINPUT4), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n333), .B1(new_n308), .B2(new_n319), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n338), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n359), .B(new_n338), .C1(new_n346), .C2(new_n354), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(new_n360), .A3(new_n363), .ZN(new_n366));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT22), .ZN(new_n368));
  INV_X1    g167(.A(G211gat), .ZN(new_n369));
  INV_X1    g168(.A(G218gat), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n372), .B2(new_n373), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n381));
  NOR2_X1   g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT25), .ZN(new_n385));
  AND2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n386), .A2(KEYINPUT24), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT69), .ZN(new_n388));
  OR2_X1    g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT69), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n386), .A2(KEYINPUT24), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT67), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n398), .A2(new_n399), .B1(KEYINPUT23), .B2(new_n382), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT68), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n387), .A2(KEYINPUT65), .A3(new_n389), .A4(new_n390), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n391), .B2(new_n393), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n402), .A2(new_n404), .A3(new_n400), .A4(new_n384), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n395), .A2(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n386), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT27), .B(G183gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT28), .ZN(new_n411));
  AOI21_X1  g210(.A(G190gat), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n382), .B(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n399), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n409), .B(new_n412), .C1(new_n410), .C2(new_n411), .ZN(new_n418));
  AND4_X1   g217(.A1(new_n408), .A2(new_n414), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT74), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n401), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT74), .ZN(new_n424));
  INV_X1    g223(.A(new_n419), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n380), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  INV_X1    g227(.A(new_n380), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n428), .A2(KEYINPUT29), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n379), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n420), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n425), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n429), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT75), .B1(new_n428), .B2(new_n380), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n433), .A2(new_n380), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n431), .B1(new_n438), .B2(new_n379), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n431), .B(new_n444), .C1(new_n438), .C2(new_n379), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(KEYINPUT30), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(KEYINPUT30), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n365), .A2(new_n366), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT31), .B(G50gat), .Z(new_n449));
  NOR3_X1   g248(.A1(new_n377), .A2(KEYINPUT29), .A3(new_n378), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n325), .B1(new_n450), .B2(KEYINPUT3), .ZN(new_n451));
  INV_X1    g250(.A(G228gat), .ZN(new_n452));
  INV_X1    g251(.A(G233gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT29), .B1(new_n319), .B2(new_n330), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n451), .B(new_n454), .C1(new_n455), .C2(new_n379), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  INV_X1    g256(.A(new_n379), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n323), .A2(new_n330), .A3(new_n324), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT29), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n454), .A4(new_n451), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n372), .A2(new_n376), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n375), .A2(new_n367), .A3(new_n371), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT29), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n325), .B1(KEYINPUT3), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n455), .B2(new_n379), .ZN(new_n467));
  INV_X1    g266(.A(new_n454), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G22gat), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n457), .A2(new_n462), .A3(new_n469), .A4(new_n204), .ZN(new_n472));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n449), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(new_n473), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n480));
  INV_X1    g279(.A(new_n449), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n448), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n485));
  NAND3_X1  g284(.A1(new_n334), .A2(new_n339), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n334), .A2(new_n339), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n340), .A2(new_n341), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT39), .B1(new_n489), .B2(new_n339), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n359), .B(new_n486), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n487), .B(KEYINPUT39), .C1(new_n339), .C2(new_n489), .ZN(new_n494));
  INV_X1    g293(.A(new_n492), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n359), .A3(new_n486), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n361), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n446), .A2(new_n447), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n362), .A2(new_n364), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n336), .B1(new_n342), .B2(KEYINPUT79), .ZN(new_n501));
  INV_X1    g300(.A(new_n353), .ZN(new_n502));
  OAI22_X1  g301(.A1(new_n352), .A2(KEYINPUT78), .B1(new_n320), .B2(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n501), .B(new_n345), .C1(new_n504), .C2(new_n347), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n359), .B1(new_n505), .B2(new_n338), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n366), .B(new_n445), .C1(new_n500), .C2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n444), .A2(KEYINPUT38), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n427), .A2(new_n430), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT37), .B1(new_n509), .B2(new_n379), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n438), .A2(new_n458), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n431), .B(new_n513), .C1(new_n438), .C2(new_n379), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n514), .B(KEYINPUT84), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n444), .B1(new_n439), .B2(KEYINPUT37), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT38), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n499), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n484), .B1(new_n524), .B2(new_n483), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n428), .A2(new_n329), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n308), .B1(new_n407), .B2(new_n419), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n529));
  NAND2_X1  g328(.A1(G227gat), .A2(G233gat), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n526), .A2(new_n527), .A3(G227gat), .A4(G233gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT32), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G15gat), .B(G43gat), .Z(new_n538));
  XNOR2_X1  g337(.A(G71gat), .B(G99gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n534), .B(KEYINPUT32), .C1(new_n536), .C2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n533), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n533), .B1(new_n543), .B2(new_n541), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT36), .B1(new_n544), .B2(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n476), .A2(new_n482), .A3(new_n546), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n553), .B(new_n448), .C1(new_n554), .C2(KEYINPUT35), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n476), .A2(new_n482), .A3(new_n546), .A4(new_n554), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n366), .B1(new_n500), .B2(new_n506), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n498), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n476), .A2(new_n482), .A3(new_n546), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n556), .B(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n295), .B1(new_n552), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  NAND2_X1  g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n570), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT94), .A3(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n568), .B1(new_n570), .B2(KEYINPUT93), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n575), .B1(KEYINPUT93), .B2(new_n568), .C1(new_n564), .C2(new_n565), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n216), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT96), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n578), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT95), .Z(new_n584));
  AND2_X1   g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n582), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n589), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n592), .B2(new_n597), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n581), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n580), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G134gat), .B(G162gat), .Z(new_n606));
  NAND2_X1  g405(.A1(G99gat), .A2(G106gat), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  INV_X1    g415(.A(G99gat), .ZN(new_n617));
  INV_X1    g416(.A(G106gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n607), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n615), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n616), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n613), .A2(new_n614), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(KEYINPUT97), .A3(new_n607), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n610), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n621), .B(new_n625), .C1(new_n240), .C2(new_n245), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n253), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n628), .A2(KEYINPUT98), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT98), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n606), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(new_n606), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n605), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n574), .A2(new_n576), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n627), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n577), .A2(new_n621), .A3(new_n625), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n650), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT100), .B1(new_n650), .B2(new_n652), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(new_n660), .A3(new_n649), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n647), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(KEYINPUT99), .A3(new_n662), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n652), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n652), .B1(new_n661), .B2(new_n662), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n658), .B1(new_n655), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n563), .A2(new_n646), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n558), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n210), .ZN(G1324gat));
  OAI21_X1  g475(.A(G8gat), .B1(new_n674), .B2(new_n498), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT16), .B(G8gat), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n674), .A2(new_n498), .A3(new_n679), .ZN(new_n680));
  MUX2_X1   g479(.A(new_n678), .B(KEYINPUT42), .S(new_n680), .Z(G1325gat));
  AND3_X1   g480(.A1(new_n548), .A2(KEYINPUT101), .A3(new_n549), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT101), .B1(new_n548), .B2(new_n549), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n674), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n546), .A2(new_n206), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n674), .B2(new_n686), .ZN(G1326gat));
  INV_X1    g486(.A(new_n483), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n674), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT43), .B(G22gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n605), .A2(new_n673), .ZN(new_n692));
  INV_X1    g491(.A(new_n645), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n563), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G29gat), .ZN(new_n696));
  INV_X1    g495(.A(new_n558), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n688), .A2(new_n559), .ZN(new_n700));
  INV_X1    g499(.A(new_n508), .ZN(new_n701));
  INV_X1    g500(.A(new_n510), .ZN(new_n702));
  INV_X1    g501(.A(new_n511), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n515), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n706), .A2(new_n365), .A3(new_n366), .A4(new_n445), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n520), .B2(new_n521), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n707), .A2(new_n709), .B1(new_n498), .B2(new_n497), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n700), .B1(new_n710), .B2(new_n688), .ZN(new_n711));
  INV_X1    g510(.A(new_n684), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n562), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n645), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n693), .B1(new_n552), .B2(new_n562), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n287), .A2(new_n293), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n287), .B2(new_n293), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n692), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n720), .A2(new_n558), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n699), .B1(new_n696), .B2(new_n727), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n498), .A2(G36gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n695), .A2(new_n729), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n730), .A2(KEYINPUT104), .A3(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n730), .B2(KEYINPUT46), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(new_n732), .B1(KEYINPUT46), .B2(new_n730), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n720), .A2(new_n498), .A3(new_n726), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  OAI21_X1  g534(.A(G36gat), .B1(new_n734), .B2(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n563), .A2(new_n220), .A3(new_n546), .A4(new_n694), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n555), .A2(new_n561), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n525), .B2(new_n684), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(new_n693), .A3(new_n714), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n562), .B1(new_n711), .B2(new_n550), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n718), .B1(new_n744), .B2(new_n645), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n712), .B(new_n725), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n738), .B1(new_n740), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n220), .B1(new_n746), .B2(KEYINPUT107), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n719), .A2(new_n751), .A3(new_n712), .A4(new_n725), .ZN(new_n752));
  AOI211_X1 g551(.A(KEYINPUT108), .B(new_n749), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(G43gat), .A3(new_n752), .ZN(new_n756));
  INV_X1    g555(.A(new_n749), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n748), .B1(new_n753), .B2(new_n758), .ZN(G1330gat));
  NOR3_X1   g558(.A1(new_n720), .A2(new_n688), .A3(new_n726), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT109), .B1(new_n760), .B2(new_n218), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n695), .A2(new_n218), .A3(new_n483), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n760), .B2(new_n218), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI221_X1 g564(.A(new_n762), .B1(KEYINPUT109), .B2(KEYINPUT48), .C1(new_n760), .C2(new_n218), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NAND3_X1  g566(.A1(new_n646), .A2(new_n672), .A3(new_n724), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n742), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  INV_X1    g569(.A(new_n768), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n713), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n697), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  INV_X1    g574(.A(new_n498), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT49), .B(G64gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT111), .ZN(G1333gat));
  NAND3_X1  g581(.A1(new_n769), .A2(new_n772), .A3(new_n546), .ZN(new_n783));
  AOI21_X1  g582(.A(G71gat), .B1(new_n783), .B2(KEYINPUT112), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT112), .B2(new_n783), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n773), .A2(G71gat), .A3(new_n712), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n483), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n742), .A2(new_n693), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n605), .A2(new_n724), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT113), .Z(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n697), .A2(new_n608), .A3(new_n672), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n672), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n720), .A2(new_n558), .A3(new_n804), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n802), .A2(new_n803), .B1(new_n805), .B2(new_n608), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n720), .A2(new_n498), .A3(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n776), .A2(new_n609), .A3(new_n672), .ZN(new_n809));
  OAI221_X1 g608(.A(new_n807), .B1(new_n808), .B2(new_n609), .C1(new_n802), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(new_n609), .ZN(new_n811));
  INV_X1    g610(.A(new_n801), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(new_n799), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n546), .A2(new_n617), .A3(new_n672), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n720), .A2(new_n684), .A3(new_n804), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n802), .A2(new_n816), .B1(new_n817), .B2(new_n617), .ZN(G1338gat));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n720), .A2(new_n688), .A3(new_n804), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n483), .A2(new_n618), .A3(new_n672), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n819), .B1(new_n820), .B2(new_n618), .C1(new_n802), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n618), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n812), .B2(new_n799), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(G1339gat));
  AND2_X1   g625(.A1(new_n602), .A2(new_n604), .ZN(new_n827));
  INV_X1    g626(.A(new_n658), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n670), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n663), .B2(new_n651), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n667), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n830), .B(KEYINPUT55), .C1(new_n667), .C2(new_n831), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n669), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n294), .A2(KEYINPUT102), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n287), .A2(new_n293), .A3(new_n721), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n291), .A2(new_n292), .A3(new_n279), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n259), .B1(new_n246), .B2(new_n256), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n841), .A2(new_n842), .B1(new_n274), .B2(new_n266), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n285), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n840), .A2(new_n672), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n840), .A2(new_n672), .A3(new_n845), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n848), .B(new_n849), .C1(new_n724), .C2(new_n836), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n850), .A3(new_n693), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n840), .A2(new_n845), .ZN(new_n852));
  INV_X1    g651(.A(new_n836), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n645), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n827), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n646), .A2(new_n673), .A3(new_n724), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n558), .A3(new_n776), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n553), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n295), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n724), .A2(G113gat), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT116), .Z(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(G1340gat));
  OAI21_X1  g663(.A(G120gat), .B1(new_n860), .B2(new_n673), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n673), .A2(G120gat), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT117), .Z(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n860), .B2(new_n867), .ZN(G1341gat));
  NOR2_X1   g667(.A1(new_n860), .A2(new_n605), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(G127gat), .Z(G1342gat));
  AOI21_X1  g669(.A(new_n560), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n859), .A2(new_n645), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n872), .B(new_n873), .Z(G1343gat));
  NAND2_X1  g673(.A1(new_n294), .A2(new_n853), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n849), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n836), .B1(new_n287), .B2(new_n293), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT118), .B1(new_n878), .B2(new_n846), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n693), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n827), .B1(new_n880), .B2(new_n854), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n856), .B1(new_n881), .B2(KEYINPUT119), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n883), .B(new_n827), .C1(new_n880), .C2(new_n854), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n483), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n886));
  INV_X1    g685(.A(new_n724), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n888), .B(new_n483), .C1(new_n855), .C2(new_n857), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n712), .A2(new_n558), .A3(new_n776), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n712), .A2(new_n688), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n295), .A2(G141gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n891), .B2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT58), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n859), .A2(new_n893), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT58), .B1(new_n899), .B2(new_n894), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n886), .A2(new_n294), .A3(new_n889), .A4(new_n890), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G141gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n898), .A2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n673), .A2(G148gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n859), .A2(new_n893), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n645), .A2(new_n853), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT123), .Z(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n852), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n827), .B1(new_n913), .B2(new_n880), .ZN(new_n914));
  NOR4_X1   g713(.A1(new_n605), .A2(new_n645), .A3(new_n294), .A4(new_n672), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n888), .B(new_n483), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n858), .B2(new_n688), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n890), .B(KEYINPUT122), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n672), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n910), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n910), .A2(G148gat), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n672), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n909), .B1(new_n920), .B2(new_n923), .ZN(G1345gat));
  AND3_X1   g723(.A1(new_n859), .A2(new_n827), .A3(new_n893), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G155gat), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n605), .A2(new_n310), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT125), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n927), .A2(new_n928), .B1(new_n922), .B2(new_n930), .ZN(G1346gat));
  NAND3_X1  g730(.A1(new_n899), .A2(new_n311), .A3(new_n645), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n922), .A2(new_n645), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n311), .ZN(G1347gat));
  INV_X1    g733(.A(new_n858), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n697), .A2(new_n498), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n553), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n283), .A3(new_n295), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n858), .A2(new_n697), .A3(new_n498), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n553), .A3(new_n887), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n940), .B2(new_n283), .ZN(G1348gat));
  NOR2_X1   g740(.A1(new_n937), .A2(new_n673), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(G176gat), .Z(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n937), .B2(new_n605), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n939), .A2(new_n409), .A3(new_n553), .A4(new_n827), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n939), .A2(new_n553), .A3(new_n645), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n948), .B2(G190gat), .ZN(new_n952));
  OAI22_X1  g751(.A1(new_n951), .A2(new_n952), .B1(G190gat), .B2(new_n948), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n893), .A3(new_n936), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n887), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n916), .A2(new_n917), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n684), .A2(new_n936), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n294), .A2(G197gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n672), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G204gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n673), .A2(G204gat), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n939), .A2(KEYINPUT126), .A3(new_n893), .A4(new_n965), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT62), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n369), .A3(new_n827), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n916), .A2(new_n917), .A3(new_n827), .A4(new_n958), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(new_n370), .B1(new_n954), .B2(new_n693), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n957), .A2(G218gat), .A3(new_n645), .A4(new_n958), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(G1355gat));
endmodule


