//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT78), .A2(G107), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT78), .A2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(G104), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT79), .A3(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G101), .B1(new_n194), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT80), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n198), .B2(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n196), .B2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n192), .A2(new_n203), .A3(G104), .A4(new_n193), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(G101), .C1(new_n194), .C2(new_n200), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n202), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  OAI211_X1 g032(.A(G128), .B(new_n215), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(new_n221), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n202), .A2(KEYINPUT82), .A3(new_n208), .A4(new_n210), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n210), .A2(new_n208), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT78), .A2(G107), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT78), .A2(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n196), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(new_n197), .A3(new_n199), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n209), .B1(new_n232), .B2(G101), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT64), .A3(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT64), .A2(G131), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n240), .A2(new_n242), .A3(new_n246), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n207), .B1(new_n205), .B2(new_n206), .ZN(new_n251));
  MUX2_X1   g065(.A(new_n250), .B(KEYINPUT4), .S(new_n251), .Z(new_n252));
  NAND4_X1  g066(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT0), .A4(G128), .ZN(new_n253));
  XNOR2_X1  g067(.A(G143), .B(G146), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT0), .B(G128), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n227), .A2(new_n237), .A3(new_n249), .A4(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(G227), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(new_n224), .C1(new_n228), .C2(new_n233), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n211), .B2(new_n224), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n235), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(KEYINPUT84), .A3(KEYINPUT12), .A4(new_n248), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n211), .A2(new_n224), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n224), .B1(new_n228), .B2(new_n233), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT83), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n275), .B2(new_n267), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n276), .B2(new_n249), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n267), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n249), .B1(new_n279), .B2(new_n235), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT84), .B1(new_n280), .B2(KEYINPUT12), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n265), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n227), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n237), .A2(new_n258), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n248), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n259), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n263), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G469), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n190), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n282), .B2(new_n287), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT85), .A3(new_n289), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n259), .B1(new_n278), .B2(new_n281), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n263), .B(KEYINPUT77), .Z(new_n297));
  AOI22_X1  g111(.A1(new_n296), .A2(new_n297), .B1(new_n265), .B2(new_n285), .ZN(new_n298));
  OAI21_X1  g112(.A(G469), .B1(new_n298), .B2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n191), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n302));
  INV_X1    g116(.A(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G116), .ZN(new_n304));
  OAI21_X1  g118(.A(G113), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G116), .B(G119), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n302), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT2), .B(G113), .Z(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n213), .A2(new_n226), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n306), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n304), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT2), .B(G113), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n252), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n310), .A2(new_n318), .A3(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT6), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n310), .B2(new_n318), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n301), .B(new_n323), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n324), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n256), .A2(G125), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n225), .B2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n332), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G210), .B1(G237), .B2(G902), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n339), .B(KEYINPUT91), .Z(new_n340));
  XNOR2_X1  g154(.A(new_n321), .B(KEYINPUT8), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n309), .A2(new_n234), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n305), .A2(KEYINPUT88), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n305), .B2(KEYINPUT88), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n311), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n211), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n343), .B1(new_n348), .B2(KEYINPUT89), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(KEYINPUT89), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n342), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n331), .A2(KEYINPUT90), .B1(KEYINPUT7), .B2(new_n335), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(new_n332), .Z(new_n353));
  NAND2_X1  g167(.A1(new_n324), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n190), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n340), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G214), .B1(G237), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n340), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n336), .B1(new_n327), .B2(new_n329), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n355), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT19), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(new_n217), .C1(new_n373), .C2(new_n370), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT16), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n364), .A3(G125), .ZN(new_n377));
  OAI211_X1 g191(.A(G146), .B(new_n377), .C1(new_n368), .C2(new_n376), .ZN(new_n378));
  NOR2_X1   g192(.A1(G237), .A2(G953), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(G143), .A3(G214), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G143), .B1(new_n379), .B2(G214), .ZN(new_n382));
  OAI21_X1  g196(.A(G131), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G214), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n214), .ZN(new_n385));
  INV_X1    g199(.A(G131), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n380), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n375), .A2(new_n378), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n369), .A2(new_n372), .A3(new_n217), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n217), .B2(new_n370), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT18), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n385), .A2(new_n380), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT18), .B(G131), .C1(new_n381), .C2(new_n382), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n196), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT17), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n383), .A2(new_n387), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT92), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n377), .B1(new_n368), .B2(new_n376), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n217), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n405), .A2(new_n378), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT92), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n383), .A2(new_n387), .A3(new_n407), .A4(new_n401), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n383), .A2(new_n401), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n403), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n398), .A3(new_n395), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n363), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT20), .B(new_n415), .C1(new_n400), .C2(new_n411), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n395), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  INV_X1    g234(.A(G475), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT93), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n424));
  OAI221_X1 g238(.A(new_n424), .B1(new_n420), .B2(new_n421), .C1(new_n414), .C2(new_n416), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT95), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT94), .A2(G122), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(KEYINPUT94), .A2(G122), .ZN(new_n430));
  OAI21_X1  g244(.A(G116), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n229), .A2(new_n230), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n312), .A2(G122), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n431), .B2(new_n433), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n427), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT13), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(G134), .C1(new_n214), .C2(G128), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G134), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n222), .A2(G143), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n214), .A2(G128), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n442), .A2(new_n443), .A3(new_n239), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n439), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n438), .A2(new_n214), .A3(G128), .A4(G134), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n430), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n312), .B1(new_n448), .B2(new_n428), .ZN(new_n449));
  INV_X1    g263(.A(new_n433), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n449), .A2(new_n450), .B1(new_n230), .B2(new_n229), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n434), .A3(KEYINPUT95), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n437), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT69), .B(G217), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n189), .A2(new_n261), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n433), .B(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(G107), .B1(new_n458), .B2(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n434), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n441), .A2(new_n444), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n431), .A2(KEYINPUT96), .A3(new_n432), .A4(new_n433), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n459), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT97), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT97), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n453), .A2(new_n457), .A3(new_n467), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n453), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n456), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n190), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT98), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(KEYINPUT98), .A3(new_n190), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n472), .A2(new_n476), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n481), .A2(G952), .A3(new_n261), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(G898), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n426), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n362), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n405), .A2(new_n378), .ZN(new_n489));
  INV_X1    g303(.A(G110), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT24), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT24), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G110), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT70), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT70), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n303), .A2(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n222), .A2(G119), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n303), .B2(G128), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n501), .A2(new_n496), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n489), .B(new_n499), .C1(new_n490), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n390), .A2(new_n378), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(KEYINPUT71), .A3(new_n490), .A4(new_n503), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n498), .B1(new_n494), .B2(new_n495), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(new_n503), .A3(new_n490), .A4(new_n496), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n506), .A2(KEYINPUT73), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT73), .B1(new_n506), .B2(new_n512), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n516), .B(new_n517), .Z(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n505), .B(new_n518), .C1(new_n513), .C2(new_n514), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n190), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n190), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n454), .B1(G234), .B2(new_n190), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n488), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT75), .B(new_n531), .C1(new_n525), .C2(new_n527), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n529), .A2(G902), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n520), .A2(new_n521), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n248), .A2(new_n257), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n240), .A2(new_n242), .A3(new_n386), .A4(new_n243), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n239), .A2(G137), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n241), .A2(G134), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n219), .A2(new_n538), .A3(new_n541), .A4(new_n223), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n311), .A2(KEYINPUT66), .A3(new_n316), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT66), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n317), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n537), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n543), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT66), .B1(new_n311), .B2(new_n316), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(KEYINPUT28), .A3(new_n537), .A4(new_n542), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n537), .A2(new_n542), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n317), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT26), .B(G101), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n379), .A2(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n546), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n256), .B1(new_n245), .B2(new_n247), .ZN(new_n563));
  INV_X1    g377(.A(new_n542), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT65), .B(KEYINPUT30), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n537), .A2(new_n542), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n562), .B1(new_n569), .B2(new_n317), .ZN(new_n570));
  INV_X1    g384(.A(new_n560), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT31), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n565), .A2(new_n568), .B1(new_n316), .B2(new_n311), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n574));
  NOR4_X1   g388(.A1(new_n573), .A2(new_n574), .A3(new_n562), .A4(new_n560), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n561), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n577), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n563), .A2(new_n564), .B1(new_n549), .B2(new_n550), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n546), .A2(new_n579), .A3(KEYINPUT68), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n553), .B(new_n581), .C1(new_n549), .C2(new_n550), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT28), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(KEYINPUT29), .A3(new_n571), .A4(new_n548), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n570), .A2(new_n571), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n555), .B2(new_n560), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n584), .B(new_n190), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n577), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n536), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n300), .A2(new_n487), .A3(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT99), .B(G101), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G3));
  INV_X1    g411(.A(new_n485), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n357), .A2(new_n361), .A3(new_n358), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n576), .A2(new_n190), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(G472), .B1(new_n576), .B2(new_n577), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n599), .A2(new_n536), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n300), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n469), .B2(new_n456), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n471), .A2(new_n606), .B1(new_n465), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(G478), .A3(new_n190), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n426), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n416), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n414), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n412), .A2(KEYINPUT100), .A3(new_n363), .A4(new_n413), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n422), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n480), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n604), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  NAND2_X1  g439(.A1(new_n528), .A2(new_n529), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT75), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n528), .A2(new_n488), .A3(new_n529), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n515), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n515), .A2(new_n630), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n534), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n300), .A2(new_n487), .A3(new_n601), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  AOI21_X1  g452(.A(new_n264), .B1(new_n285), .B2(new_n259), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n270), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT84), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n277), .A3(new_n271), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n639), .B1(new_n643), .B2(new_n265), .ZN(new_n644));
  NOR4_X1   g458(.A1(new_n644), .A2(new_n291), .A3(G469), .A4(G902), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT85), .B1(new_n293), .B2(new_n289), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n299), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n191), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n578), .A2(new_n589), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n592), .A2(new_n591), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n533), .A2(new_n634), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n647), .A2(new_n648), .A3(new_n362), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n482), .B1(new_n483), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n621), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n222), .ZN(G30));
  AOI21_X1  g472(.A(new_n340), .B1(new_n338), .B2(new_n356), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n360), .A2(new_n359), .A3(new_n355), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT38), .ZN(new_n662));
  INV_X1    g476(.A(new_n358), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n478), .B2(new_n479), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n426), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT103), .B1(new_n635), .B2(new_n665), .ZN(new_n666));
  OR3_X1    g480(.A1(new_n635), .A2(new_n665), .A3(KEYINPUT103), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n662), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n570), .A2(new_n571), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n580), .A2(new_n582), .A3(new_n560), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n190), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n650), .A2(new_n673), .A3(new_n578), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n592), .A2(new_n591), .B1(G472), .B2(new_n672), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT101), .B1(new_n677), .B2(new_n578), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n654), .B(KEYINPUT39), .Z(new_n681));
  AND3_X1   g495(.A1(new_n647), .A2(new_n648), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n668), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n674), .B(new_n675), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT102), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n662), .A2(new_n667), .A3(new_n666), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  INV_X1    g506(.A(new_n686), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n692), .A3(new_n693), .A4(new_n684), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n214), .ZN(G45));
  INV_X1    g510(.A(new_n654), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n426), .A2(new_n610), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n652), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n217), .ZN(G48));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n644), .B2(G902), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n293), .A2(KEYINPUT105), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(G469), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n295), .A2(new_n648), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n295), .A2(KEYINPUT106), .A3(new_n704), .A4(new_n648), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n599), .A2(new_n611), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n594), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NOR2_X1   g526(.A1(new_n599), .A2(new_n621), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n594), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n648), .A2(new_n295), .A3(new_n362), .A4(new_n704), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n651), .A2(new_n486), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n295), .A2(new_n362), .A3(new_n648), .A4(new_n704), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n718), .A3(KEYINPUT107), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n303), .ZN(G21));
  AND2_X1   g538(.A1(new_n583), .A2(new_n548), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n725), .A2(new_n571), .B1(new_n572), .B2(new_n575), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n600), .A2(G472), .B1(new_n577), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n533), .A2(new_n535), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n357), .A2(new_n361), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n728), .A2(new_n729), .A3(new_n665), .A4(new_n485), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n707), .A2(new_n708), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n635), .A2(new_n727), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n698), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n717), .A2(KEYINPUT108), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  INV_X1    g550(.A(new_n698), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n635), .A3(new_n727), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n721), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n650), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT111), .B1(new_n592), .B2(new_n591), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n590), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n536), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT112), .B1(new_n745), .B2(new_n536), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n647), .A2(KEYINPUT109), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(new_n299), .C1(new_n645), .C2(new_n646), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n648), .A2(new_n358), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n661), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n751), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n752), .A2(new_n594), .A3(new_n754), .A4(new_n757), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n698), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  OR2_X1    g578(.A1(new_n761), .A2(new_n656), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NAND3_X1  g580(.A1(new_n610), .A2(new_n425), .A3(new_n423), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT43), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n602), .A3(new_n635), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n358), .B1(new_n659), .B2(new_n660), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n778));
  OAI21_X1  g592(.A(G469), .B1(new_n298), .B2(KEYINPUT45), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n298), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n778), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n784), .A2(KEYINPUT114), .A3(KEYINPUT46), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n295), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n777), .A2(new_n791), .A3(new_n648), .A4(new_n681), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n648), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(KEYINPUT47), .A3(new_n648), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n776), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n593), .A2(new_n799), .A3(new_n536), .A4(new_n737), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NOR4_X1   g616(.A1(new_n662), .A2(new_n767), .A3(new_n536), .A4(new_n756), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n295), .A2(new_n704), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT49), .Z(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n805), .A3(new_n689), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n710), .B(new_n714), .C1(new_n720), .C2(new_n722), .ZN(new_n807));
  INV_X1    g621(.A(new_n480), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n611), .B1(new_n426), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n300), .A2(new_n603), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n731), .A2(new_n595), .A3(new_n636), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n808), .A2(new_n620), .A3(new_n697), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n776), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n808), .A2(new_n620), .A3(new_n697), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n358), .A4(new_n729), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n300), .A2(new_n815), .A3(new_n817), .A4(new_n651), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n752), .A2(new_n734), .A3(new_n754), .A4(new_n757), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n818), .B(new_n819), .C1(new_n761), .C2(new_n656), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n762), .B2(new_n759), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n191), .A2(new_n654), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n357), .A2(new_n361), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n635), .A3(new_n665), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n752), .A2(new_n688), .A3(new_n754), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n426), .A2(new_n664), .ZN(new_n830));
  INV_X1    g644(.A(new_n634), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n530), .A2(new_n532), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n661), .A2(new_n830), .A3(new_n832), .A4(new_n824), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n679), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(KEYINPUT116), .A3(new_n752), .A4(new_n754), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n652), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n655), .B2(new_n737), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n740), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n823), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n652), .B1(new_n656), .B2(new_n698), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n739), .B2(new_n735), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n822), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT52), .A2(new_n836), .A3(new_n740), .A4(new_n839), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n843), .B2(new_n836), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n821), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n841), .A2(new_n854), .A3(new_n844), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n848), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n846), .A2(new_n847), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n855), .A3(new_n822), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n859), .B2(new_n847), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n860), .B2(new_n849), .ZN(new_n861));
  INV_X1    g675(.A(new_n482), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n770), .A2(new_n862), .A3(new_n728), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n804), .A2(new_n648), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n799), .B(new_n863), .C1(new_n798), .C2(new_n864), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n804), .A2(new_n661), .A3(new_n862), .A4(new_n756), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n771), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n733), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n689), .A2(new_n866), .A3(new_n747), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n426), .A2(new_n610), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n662), .A2(new_n358), .ZN(new_n873));
  INV_X1    g687(.A(new_n804), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n648), .A3(new_n874), .A4(new_n863), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT50), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT51), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n866), .A2(new_n751), .A3(new_n771), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n869), .A2(new_n612), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n261), .A2(G952), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n863), .B2(new_n717), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI211_X1 g702(.A(KEYINPUT120), .B(KEYINPUT48), .C1(new_n881), .C2(new_n882), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n865), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n877), .A2(KEYINPUT118), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n872), .B2(new_n876), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT51), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n890), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n861), .A2(new_n878), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n806), .B1(new_n897), .B2(new_n898), .ZN(G75));
  NOR2_X1   g713(.A1(new_n261), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n190), .B1(new_n848), .B2(new_n856), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(new_n340), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n330), .B(new_n337), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n901), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n903), .B2(new_n906), .ZN(G51));
  AOI211_X1 g722(.A(new_n190), .B(new_n784), .C1(new_n848), .C2(new_n856), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n288), .B(KEYINPUT121), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n852), .A2(new_n855), .A3(new_n853), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n822), .B2(new_n845), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n857), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n785), .B(KEYINPUT57), .Z(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n909), .B1(new_n916), .B2(KEYINPUT122), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n918));
  INV_X1    g732(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n913), .B2(new_n857), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n900), .B1(new_n917), .B2(new_n921), .ZN(G54));
  AND2_X1   g736(.A1(KEYINPUT58), .A2(G475), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n902), .A2(new_n412), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n412), .B1(new_n902), .B2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n900), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT59), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n608), .B1(new_n861), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n914), .A2(new_n608), .A3(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n900), .ZN(G63));
  NAND2_X1  g745(.A1(new_n848), .A2(new_n856), .ZN(new_n932));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n633), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n901), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n520), .A2(new_n521), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT123), .Z(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n932), .B2(new_n934), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n936), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(G953), .B1(new_n484), .B2(new_n333), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n812), .B2(G953), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n327), .B(new_n329), .C1(G898), .C2(new_n261), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  AOI211_X1 g761(.A(new_n729), .B(new_n665), .C1(new_n749), .C2(new_n750), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n791), .A2(new_n648), .A3(new_n681), .A4(new_n948), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n763), .A2(new_n949), .A3(new_n765), .A4(new_n843), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n801), .A2(new_n950), .A3(new_n261), .A4(new_n792), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n374), .B1(new_n373), .B2(new_n370), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n569), .B(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(G900), .B2(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n809), .B(KEYINPUT125), .Z(new_n958));
  AND4_X1   g772(.A1(new_n594), .A2(new_n958), .A3(new_n682), .A4(new_n799), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n695), .B2(new_n840), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n687), .A2(new_n694), .A3(KEYINPUT62), .A4(new_n843), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n792), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n798), .B2(new_n800), .ZN(new_n965));
  AOI21_X1  g779(.A(G953), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n953), .B(KEYINPUT124), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n955), .B(new_n957), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n955), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n972), .A2(KEYINPUT127), .A3(new_n956), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT127), .B1(new_n972), .B2(new_n956), .ZN(new_n974));
  OAI22_X1  g788(.A1(new_n970), .A2(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G72));
  INV_X1    g789(.A(new_n585), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n669), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n965), .A2(new_n950), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n560), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n963), .A2(new_n965), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(new_n812), .C1(new_n980), .C2(new_n560), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  AOI21_X1  g797(.A(new_n977), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n983), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n901), .B1(new_n860), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(G57));
endmodule


